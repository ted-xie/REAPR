library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Brill is
	port (
		clock, reset, run : in std_logic;
		data_in : in std_logic_vector(7 downto 0);
		reports : out std_logic_vector(218-1 downto 0)
	);
end Brill;

architecture Structure of Brill is
	--------------------------
	-- Component Declarations
	--------------------------
	COMPONENT ste_sim
		PORT
		(
			bitvector	:	in std_logic_vector(255 downto 0);
			char_in		:	in std_logic_vector(7 downto 0);
			clock, reset, run		:	in std_logic;
			Enable	:	in std_logic;
			match		:	out std_logic
		);
	END COMPONENT;
	COMPONENT Counter
		GENERIC	(target : INTEGER := 8;
			at_target : INTEGER := 0);
		PORT	(clock : IN std_logic;
			Enable, Reset, run : IN std_logic;
--			q : OUT std_logic_vector(11 DOWNTO 0);
			match : OUT std_logic);
	END COMPONENT;
	--------------------------
	-- Signal Declarations
	--------------------------
	--- STEs
	signal bitvectord2d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2d : std_logic := '1';
	signal matchd2d : std_logic := '0';
	
	signal bitvectord3d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3d : std_logic := '0';
	signal matchd3d : std_logic := '0';
	
	signal bitvectord4d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled4d : std_logic := '0';
	signal matchd4d : std_logic := '0';
	
	signal bitvectord5d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled5d : std_logic := '0';
	signal matchd5d : std_logic := '0';
	
	signal bitvectord6d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled6d : std_logic := '0';
	signal matchd6d : std_logic := '0';
	
	signal bitvectord7d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled7d : std_logic := '0';
	signal matchd7d : std_logic := '0';
	
	signal bitvectord8d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled8d : std_logic := '0';
	signal matchd8d : std_logic := '0';
	
	signal bitvectord9d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled9d : std_logic := '0';
	signal matchd9d : std_logic := '0';
	
	signal bitvectord10d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled10d : std_logic := '0';
	signal matchd10d : std_logic := '0';
	
	signal bitvectord11d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled11d : std_logic := '0';
	signal matchd11d : std_logic := '0';
	
	signal bitvectord12d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled12d : std_logic := '0';
	signal matchd12d : std_logic := '0';
	
	signal bitvectord13d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled13d : std_logic := '0';
	signal matchd13d : std_logic := '0';
	
	signal bitvectord14d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled14d : std_logic := '0';
	signal matchd14d : std_logic := '0';
	
	signal bitvectord15d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled15d : std_logic := '0';
	signal matchd15d : std_logic := '0';
	
	signal bitvectord16d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled16d : std_logic := '0';
	signal matchd16d : std_logic := '0';
	
	signal bitvectord17d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled17d : std_logic := '1';
	signal matchd17d : std_logic := '0';
	
	signal bitvectord18d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled18d : std_logic := '0';
	signal matchd18d : std_logic := '0';
	
	signal bitvectord19d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled19d : std_logic := '0';
	signal matchd19d : std_logic := '0';
	
	signal bitvectord20d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled20d : std_logic := '0';
	signal matchd20d : std_logic := '0';
	
	signal bitvectord21d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled21d : std_logic := '0';
	signal matchd21d : std_logic := '0';
	
	signal bitvectord22d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled22d : std_logic := '0';
	signal matchd22d : std_logic := '0';
	
	signal bitvectord23d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled23d : std_logic := '0';
	signal matchd23d : std_logic := '0';
	
	signal bitvectord24d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled24d : std_logic := '0';
	signal matchd24d : std_logic := '0';
	
	signal bitvectord25d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled25d : std_logic := '0';
	signal matchd25d : std_logic := '0';
	
	signal bitvectord26d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled26d : std_logic := '0';
	signal matchd26d : std_logic := '0';
	
	signal bitvectord27d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled27d : std_logic := '0';
	signal matchd27d : std_logic := '0';
	
	signal bitvectord28d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled28d : std_logic := '0';
	signal matchd28d : std_logic := '0';
	
	signal bitvectord29d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled29d : std_logic := '0';
	signal matchd29d : std_logic := '0';
	
	signal bitvectord30d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled30d : std_logic := '0';
	signal matchd30d : std_logic := '0';
	
	signal bitvectord31d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled31d : std_logic := '0';
	signal matchd31d : std_logic := '0';
	
	signal bitvectord32d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled32d : std_logic := '1';
	signal matchd32d : std_logic := '0';
	
	signal bitvectord33d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled33d : std_logic := '0';
	signal matchd33d : std_logic := '0';
	
	signal bitvectord34d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled34d : std_logic := '0';
	signal matchd34d : std_logic := '0';
	
	signal bitvectord35d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled35d : std_logic := '0';
	signal matchd35d : std_logic := '0';
	
	signal bitvectord36d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled36d : std_logic := '0';
	signal matchd36d : std_logic := '0';
	
	signal bitvectord37d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled37d : std_logic := '0';
	signal matchd37d : std_logic := '0';
	
	signal bitvectord38d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled38d : std_logic := '0';
	signal matchd38d : std_logic := '0';
	
	signal bitvectord39d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled39d : std_logic := '0';
	signal matchd39d : std_logic := '0';
	
	signal bitvectord40d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled40d : std_logic := '0';
	signal matchd40d : std_logic := '0';
	
	signal bitvectord41d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled41d : std_logic := '0';
	signal matchd41d : std_logic := '0';
	
	signal bitvectord42d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled42d : std_logic := '0';
	signal matchd42d : std_logic := '0';
	
	signal bitvectord43d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled43d : std_logic := '0';
	signal matchd43d : std_logic := '0';
	
	signal bitvectord44d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled44d : std_logic := '0';
	signal matchd44d : std_logic := '0';
	
	signal bitvectord45d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled45d : std_logic := '0';
	signal matchd45d : std_logic := '0';
	
	signal bitvectord46d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled46d : std_logic := '0';
	signal matchd46d : std_logic := '0';
	
	signal bitvectord47d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled47d : std_logic := '1';
	signal matchd47d : std_logic := '0';
	
	signal bitvectord48d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000";
	signal Enabled48d : std_logic := '0';
	signal matchd48d : std_logic := '0';
	
	signal bitvectord49d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled49d : std_logic := '0';
	signal matchd49d : std_logic := '0';
	
	signal bitvectord50d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled50d : std_logic := '0';
	signal matchd50d : std_logic := '0';
	
	signal bitvectord51d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled51d : std_logic := '0';
	signal matchd51d : std_logic := '0';
	
	signal bitvectord52d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled52d : std_logic := '0';
	signal matchd52d : std_logic := '0';
	
	signal bitvectord53d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled53d : std_logic := '0';
	signal matchd53d : std_logic := '0';
	
	signal bitvectord54d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled54d : std_logic := '0';
	signal matchd54d : std_logic := '0';
	
	signal bitvectord55d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled55d : std_logic := '0';
	signal matchd55d : std_logic := '0';
	
	signal bitvectord56d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled56d : std_logic := '0';
	signal matchd56d : std_logic := '0';
	
	signal bitvectord57d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled57d : std_logic := '0';
	signal matchd57d : std_logic := '0';
	
	signal bitvectord58d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled58d : std_logic := '0';
	signal matchd58d : std_logic := '0';
	
	signal bitvectord59d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled59d : std_logic := '0';
	signal matchd59d : std_logic := '0';
	
	signal bitvectord60d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled60d : std_logic := '1';
	signal matchd60d : std_logic := '0';
	
	signal bitvectord61d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled61d : std_logic := '0';
	signal matchd61d : std_logic := '0';
	
	signal bitvectord62d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled62d : std_logic := '0';
	signal matchd62d : std_logic := '0';
	
	signal bitvectord63d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled63d : std_logic := '0';
	signal matchd63d : std_logic := '0';
	
	signal bitvectord64d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled64d : std_logic := '0';
	signal matchd64d : std_logic := '0';
	
	signal bitvectord65d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled65d : std_logic := '0';
	signal matchd65d : std_logic := '0';
	
	signal bitvectord66d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled66d : std_logic := '0';
	signal matchd66d : std_logic := '0';
	
	signal bitvectord67d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled67d : std_logic := '0';
	signal matchd67d : std_logic := '0';
	
	signal bitvectord68d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled68d : std_logic := '0';
	signal matchd68d : std_logic := '0';
	
	signal bitvectord69d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled69d : std_logic := '0';
	signal matchd69d : std_logic := '0';
	
	signal bitvectord70d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled70d : std_logic := '0';
	signal matchd70d : std_logic := '0';
	
	signal bitvectord71d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled71d : std_logic := '0';
	signal matchd71d : std_logic := '0';
	
	signal bitvectord72d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled72d : std_logic := '1';
	signal matchd72d : std_logic := '0';
	
	signal bitvectord73d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled73d : std_logic := '0';
	signal matchd73d : std_logic := '0';
	
	signal bitvectord74d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled74d : std_logic := '0';
	signal matchd74d : std_logic := '0';
	
	signal bitvectord75d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled75d : std_logic := '0';
	signal matchd75d : std_logic := '0';
	
	signal bitvectord76d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled76d : std_logic := '0';
	signal matchd76d : std_logic := '0';
	
	signal bitvectord77d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled77d : std_logic := '0';
	signal matchd77d : std_logic := '0';
	
	signal bitvectord78d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled78d : std_logic := '0';
	signal matchd78d : std_logic := '0';
	
	signal bitvectord79d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled79d : std_logic := '0';
	signal matchd79d : std_logic := '0';
	
	signal bitvectord80d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000";
	signal Enabled80d : std_logic := '0';
	signal matchd80d : std_logic := '0';
	
	signal bitvectord81d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled81d : std_logic := '0';
	signal matchd81d : std_logic := '0';
	
	signal bitvectord82d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000";
	signal Enabled82d : std_logic := '0';
	signal matchd82d : std_logic := '0';
	
	signal bitvectord83d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled83d : std_logic := '0';
	signal matchd83d : std_logic := '0';
	
	signal bitvectord84d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled84d : std_logic := '0';
	signal matchd84d : std_logic := '0';
	
	signal bitvectord85d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled85d : std_logic := '0';
	signal matchd85d : std_logic := '0';
	
	signal bitvectord86d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled86d : std_logic := '1';
	signal matchd86d : std_logic := '0';
	
	signal bitvectord87d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled87d : std_logic := '0';
	signal matchd87d : std_logic := '0';
	
	signal bitvectord88d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled88d : std_logic := '0';
	signal matchd88d : std_logic := '0';
	
	signal bitvectord89d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled89d : std_logic := '0';
	signal matchd89d : std_logic := '0';
	
	signal bitvectord90d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled90d : std_logic := '0';
	signal matchd90d : std_logic := '0';
	
	signal bitvectord91d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled91d : std_logic := '0';
	signal matchd91d : std_logic := '0';
	
	signal bitvectord92d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled92d : std_logic := '0';
	signal matchd92d : std_logic := '0';
	
	signal bitvectord93d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled93d : std_logic := '0';
	signal matchd93d : std_logic := '0';
	
	signal bitvectord94d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled94d : std_logic := '0';
	signal matchd94d : std_logic := '0';
	
	signal bitvectord95d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled95d : std_logic := '0';
	signal matchd95d : std_logic := '0';
	
	signal bitvectord96d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled96d : std_logic := '0';
	signal matchd96d : std_logic := '0';
	
	signal bitvectord97d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled97d : std_logic := '0';
	signal matchd97d : std_logic := '0';
	
	signal bitvectord98d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled98d : std_logic := '0';
	signal matchd98d : std_logic := '0';
	
	signal bitvectord99d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled99d : std_logic := '0';
	signal matchd99d : std_logic := '0';
	
	signal bitvectord100d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled100d : std_logic := '1';
	signal matchd100d : std_logic := '0';
	
	signal bitvectord101d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled101d : std_logic := '0';
	signal matchd101d : std_logic := '0';
	
	signal bitvectord102d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled102d : std_logic := '0';
	signal matchd102d : std_logic := '0';
	
	signal bitvectord103d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled103d : std_logic := '0';
	signal matchd103d : std_logic := '0';
	
	signal bitvectord104d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled104d : std_logic := '0';
	signal matchd104d : std_logic := '0';
	
	signal bitvectord105d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled105d : std_logic := '0';
	signal matchd105d : std_logic := '0';
	
	signal bitvectord106d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000";
	signal Enabled106d : std_logic := '0';
	signal matchd106d : std_logic := '0';
	
	signal bitvectord107d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled107d : std_logic := '0';
	signal matchd107d : std_logic := '0';
	
	signal bitvectord108d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled108d : std_logic := '0';
	signal matchd108d : std_logic := '0';
	
	signal bitvectord109d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled109d : std_logic := '0';
	signal matchd109d : std_logic := '0';
	
	signal bitvectord110d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled110d : std_logic := '0';
	signal matchd110d : std_logic := '0';
	
	signal bitvectord111d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled111d : std_logic := '1';
	signal matchd111d : std_logic := '0';
	
	signal bitvectord112d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled112d : std_logic := '0';
	signal matchd112d : std_logic := '0';
	
	signal bitvectord113d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled113d : std_logic := '0';
	signal matchd113d : std_logic := '0';
	
	signal bitvectord114d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled114d : std_logic := '0';
	signal matchd114d : std_logic := '0';
	
	signal bitvectord115d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled115d : std_logic := '0';
	signal matchd115d : std_logic := '0';
	
	signal bitvectord116d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled116d : std_logic := '0';
	signal matchd116d : std_logic := '0';
	
	signal bitvectord117d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled117d : std_logic := '0';
	signal matchd117d : std_logic := '0';
	
	signal bitvectord118d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled118d : std_logic := '0';
	signal matchd118d : std_logic := '0';
	
	signal bitvectord119d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled119d : std_logic := '0';
	signal matchd119d : std_logic := '0';
	
	signal bitvectord120d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled120d : std_logic := '0';
	signal matchd120d : std_logic := '0';
	
	signal bitvectord121d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled121d : std_logic := '0';
	signal matchd121d : std_logic := '0';
	
	signal bitvectord122d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled122d : std_logic := '0';
	signal matchd122d : std_logic := '0';
	
	signal bitvectord123d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled123d : std_logic := '1';
	signal matchd123d : std_logic := '0';
	
	signal bitvectord124d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled124d : std_logic := '0';
	signal matchd124d : std_logic := '0';
	
	signal bitvectord125d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled125d : std_logic := '0';
	signal matchd125d : std_logic := '0';
	
	signal bitvectord126d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled126d : std_logic := '0';
	signal matchd126d : std_logic := '0';
	
	signal bitvectord127d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled127d : std_logic := '0';
	signal matchd127d : std_logic := '0';
	
	signal bitvectord128d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled128d : std_logic := '0';
	signal matchd128d : std_logic := '0';
	
	signal bitvectord129d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled129d : std_logic := '0';
	signal matchd129d : std_logic := '0';
	
	signal bitvectord130d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled130d : std_logic := '0';
	signal matchd130d : std_logic := '0';
	
	signal bitvectord131d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled131d : std_logic := '0';
	signal matchd131d : std_logic := '0';
	
	signal bitvectord132d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled132d : std_logic := '0';
	signal matchd132d : std_logic := '0';
	
	signal bitvectord133d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled133d : std_logic := '0';
	signal matchd133d : std_logic := '0';
	
	signal bitvectord134d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled134d : std_logic := '0';
	signal matchd134d : std_logic := '0';
	
	signal bitvectord135d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled135d : std_logic := '0';
	signal matchd135d : std_logic := '0';
	
	signal bitvectord136d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled136d : std_logic := '0';
	signal matchd136d : std_logic := '0';
	
	signal bitvectord137d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled137d : std_logic := '0';
	signal matchd137d : std_logic := '0';
	
	signal bitvectord138d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled138d : std_logic := '1';
	signal matchd138d : std_logic := '0';
	
	signal bitvectord139d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled139d : std_logic := '0';
	signal matchd139d : std_logic := '0';
	
	signal bitvectord140d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled140d : std_logic := '0';
	signal matchd140d : std_logic := '0';
	
	signal bitvectord141d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled141d : std_logic := '0';
	signal matchd141d : std_logic := '0';
	
	signal bitvectord142d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled142d : std_logic := '0';
	signal matchd142d : std_logic := '0';
	
	signal bitvectord143d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled143d : std_logic := '0';
	signal matchd143d : std_logic := '0';
	
	signal bitvectord144d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled144d : std_logic := '0';
	signal matchd144d : std_logic := '0';
	
	signal bitvectord145d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled145d : std_logic := '0';
	signal matchd145d : std_logic := '0';
	
	signal bitvectord146d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled146d : std_logic := '0';
	signal matchd146d : std_logic := '0';
	
	signal bitvectord147d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled147d : std_logic := '0';
	signal matchd147d : std_logic := '0';
	
	signal bitvectord148d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled148d : std_logic := '0';
	signal matchd148d : std_logic := '0';
	
	signal bitvectord149d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled149d : std_logic := '0';
	signal matchd149d : std_logic := '0';
	
	signal bitvectord150d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled150d : std_logic := '0';
	signal matchd150d : std_logic := '0';
	
	signal bitvectord151d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled151d : std_logic := '0';
	signal matchd151d : std_logic := '0';
	
	signal bitvectord152d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled152d : std_logic := '1';
	signal matchd152d : std_logic := '0';
	
	signal bitvectord153d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled153d : std_logic := '0';
	signal matchd153d : std_logic := '0';
	
	signal bitvectord154d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled154d : std_logic := '0';
	signal matchd154d : std_logic := '0';
	
	signal bitvectord155d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled155d : std_logic := '0';
	signal matchd155d : std_logic := '0';
	
	signal bitvectord156d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled156d : std_logic := '0';
	signal matchd156d : std_logic := '0';
	
	signal bitvectord157d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled157d : std_logic := '0';
	signal matchd157d : std_logic := '0';
	
	signal bitvectord158d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled158d : std_logic := '0';
	signal matchd158d : std_logic := '0';
	
	signal bitvectord159d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled159d : std_logic := '0';
	signal matchd159d : std_logic := '0';
	
	signal bitvectord160d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled160d : std_logic := '0';
	signal matchd160d : std_logic := '0';
	
	signal bitvectord161d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled161d : std_logic := '0';
	signal matchd161d : std_logic := '0';
	
	signal bitvectord162d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled162d : std_logic := '0';
	signal matchd162d : std_logic := '0';
	
	signal bitvectord163d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled163d : std_logic := '0';
	signal matchd163d : std_logic := '0';
	
	signal bitvectord164d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled164d : std_logic := '0';
	signal matchd164d : std_logic := '0';
	
	signal bitvectord165d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled165d : std_logic := '0';
	signal matchd165d : std_logic := '0';
	
	signal bitvectord166d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled166d : std_logic := '1';
	signal matchd166d : std_logic := '0';
	
	signal bitvectord167d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled167d : std_logic := '0';
	signal matchd167d : std_logic := '0';
	
	signal bitvectord168d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled168d : std_logic := '0';
	signal matchd168d : std_logic := '0';
	
	signal bitvectord169d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled169d : std_logic := '0';
	signal matchd169d : std_logic := '0';
	
	signal bitvectord170d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled170d : std_logic := '0';
	signal matchd170d : std_logic := '0';
	
	signal bitvectord171d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled171d : std_logic := '0';
	signal matchd171d : std_logic := '0';
	
	signal bitvectord172d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled172d : std_logic := '0';
	signal matchd172d : std_logic := '0';
	
	signal bitvectord173d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled173d : std_logic := '0';
	signal matchd173d : std_logic := '0';
	
	signal bitvectord174d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled174d : std_logic := '0';
	signal matchd174d : std_logic := '0';
	
	signal bitvectord175d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled175d : std_logic := '0';
	signal matchd175d : std_logic := '0';
	
	signal bitvectord176d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled176d : std_logic := '0';
	signal matchd176d : std_logic := '0';
	
	signal bitvectord177d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled177d : std_logic := '1';
	signal matchd177d : std_logic := '0';
	
	signal bitvectord178d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled178d : std_logic := '0';
	signal matchd178d : std_logic := '0';
	
	signal bitvectord179d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled179d : std_logic := '0';
	signal matchd179d : std_logic := '0';
	
	signal bitvectord180d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled180d : std_logic := '0';
	signal matchd180d : std_logic := '0';
	
	signal bitvectord181d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled181d : std_logic := '0';
	signal matchd181d : std_logic := '0';
	
	signal bitvectord182d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled182d : std_logic := '0';
	signal matchd182d : std_logic := '0';
	
	signal bitvectord183d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled183d : std_logic := '0';
	signal matchd183d : std_logic := '0';
	
	signal bitvectord184d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled184d : std_logic := '0';
	signal matchd184d : std_logic := '0';
	
	signal bitvectord185d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled185d : std_logic := '0';
	signal matchd185d : std_logic := '0';
	
	signal bitvectord186d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled186d : std_logic := '0';
	signal matchd186d : std_logic := '0';
	
	signal bitvectord187d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled187d : std_logic := '0';
	signal matchd187d : std_logic := '0';
	
	signal bitvectord188d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled188d : std_logic := '1';
	signal matchd188d : std_logic := '0';
	
	signal bitvectord189d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled189d : std_logic := '0';
	signal matchd189d : std_logic := '0';
	
	signal bitvectord190d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled190d : std_logic := '0';
	signal matchd190d : std_logic := '0';
	
	signal bitvectord191d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled191d : std_logic := '0';
	signal matchd191d : std_logic := '0';
	
	signal bitvectord192d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled192d : std_logic := '0';
	signal matchd192d : std_logic := '0';
	
	signal bitvectord193d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled193d : std_logic := '0';
	signal matchd193d : std_logic := '0';
	
	signal bitvectord194d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled194d : std_logic := '0';
	signal matchd194d : std_logic := '0';
	
	signal bitvectord195d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled195d : std_logic := '0';
	signal matchd195d : std_logic := '0';
	
	signal bitvectord196d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000";
	signal Enabled196d : std_logic := '0';
	signal matchd196d : std_logic := '0';
	
	signal bitvectord197d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled197d : std_logic := '0';
	signal matchd197d : std_logic := '0';
	
	signal bitvectord198d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled198d : std_logic := '0';
	signal matchd198d : std_logic := '0';
	
	signal bitvectord199d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled199d : std_logic := '0';
	signal matchd199d : std_logic := '0';
	
	signal bitvectord200d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled200d : std_logic := '0';
	signal matchd200d : std_logic := '0';
	
	signal bitvectord201d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled201d : std_logic := '1';
	signal matchd201d : std_logic := '0';
	
	signal bitvectord202d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled202d : std_logic := '0';
	signal matchd202d : std_logic := '0';
	
	signal bitvectord203d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled203d : std_logic := '0';
	signal matchd203d : std_logic := '0';
	
	signal bitvectord204d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled204d : std_logic := '0';
	signal matchd204d : std_logic := '0';
	
	signal bitvectord205d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled205d : std_logic := '0';
	signal matchd205d : std_logic := '0';
	
	signal bitvectord206d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled206d : std_logic := '0';
	signal matchd206d : std_logic := '0';
	
	signal bitvectord207d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled207d : std_logic := '0';
	signal matchd207d : std_logic := '0';
	
	signal bitvectord208d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000";
	signal Enabled208d : std_logic := '0';
	signal matchd208d : std_logic := '0';
	
	signal bitvectord209d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled209d : std_logic := '0';
	signal matchd209d : std_logic := '0';
	
	signal bitvectord210d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled210d : std_logic := '0';
	signal matchd210d : std_logic := '0';
	
	signal bitvectord211d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled211d : std_logic := '0';
	signal matchd211d : std_logic := '0';
	
	signal bitvectord212d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled212d : std_logic := '1';
	signal matchd212d : std_logic := '0';
	
	signal bitvectord213d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled213d : std_logic := '0';
	signal matchd213d : std_logic := '0';
	
	signal bitvectord214d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled214d : std_logic := '0';
	signal matchd214d : std_logic := '0';
	
	signal bitvectord215d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled215d : std_logic := '0';
	signal matchd215d : std_logic := '0';
	
	signal bitvectord216d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled216d : std_logic := '0';
	signal matchd216d : std_logic := '0';
	
	signal bitvectord217d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled217d : std_logic := '0';
	signal matchd217d : std_logic := '0';
	
	signal bitvectord218d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled218d : std_logic := '0';
	signal matchd218d : std_logic := '0';
	
	signal bitvectord219d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled219d : std_logic := '0';
	signal matchd219d : std_logic := '0';
	
	signal bitvectord220d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled220d : std_logic := '0';
	signal matchd220d : std_logic := '0';
	
	signal bitvectord221d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled221d : std_logic := '0';
	signal matchd221d : std_logic := '0';
	
	signal bitvectord222d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled222d : std_logic := '0';
	signal matchd222d : std_logic := '0';
	
	signal bitvectord223d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled223d : std_logic := '1';
	signal matchd223d : std_logic := '0';
	
	signal bitvectord224d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled224d : std_logic := '0';
	signal matchd224d : std_logic := '0';
	
	signal bitvectord225d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled225d : std_logic := '0';
	signal matchd225d : std_logic := '0';
	
	signal bitvectord226d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled226d : std_logic := '0';
	signal matchd226d : std_logic := '0';
	
	signal bitvectord227d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled227d : std_logic := '0';
	signal matchd227d : std_logic := '0';
	
	signal bitvectord228d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled228d : std_logic := '0';
	signal matchd228d : std_logic := '0';
	
	signal bitvectord229d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled229d : std_logic := '0';
	signal matchd229d : std_logic := '0';
	
	signal bitvectord230d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled230d : std_logic := '0';
	signal matchd230d : std_logic := '0';
	
	signal bitvectord231d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled231d : std_logic := '0';
	signal matchd231d : std_logic := '0';
	
	signal bitvectord232d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled232d : std_logic := '0';
	signal matchd232d : std_logic := '0';
	
	signal bitvectord233d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled233d : std_logic := '0';
	signal matchd233d : std_logic := '0';
	
	signal bitvectord234d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled234d : std_logic := '0';
	signal matchd234d : std_logic := '0';
	
	signal bitvectord235d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled235d : std_logic := '1';
	signal matchd235d : std_logic := '0';
	
	signal bitvectord236d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled236d : std_logic := '0';
	signal matchd236d : std_logic := '0';
	
	signal bitvectord237d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled237d : std_logic := '0';
	signal matchd237d : std_logic := '0';
	
	signal bitvectord238d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled238d : std_logic := '0';
	signal matchd238d : std_logic := '0';
	
	signal bitvectord239d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled239d : std_logic := '0';
	signal matchd239d : std_logic := '0';
	
	signal bitvectord240d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled240d : std_logic := '0';
	signal matchd240d : std_logic := '0';
	
	signal bitvectord241d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled241d : std_logic := '0';
	signal matchd241d : std_logic := '0';
	
	signal bitvectord242d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled242d : std_logic := '0';
	signal matchd242d : std_logic := '0';
	
	signal bitvectord243d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled243d : std_logic := '0';
	signal matchd243d : std_logic := '0';
	
	signal bitvectord244d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled244d : std_logic := '0';
	signal matchd244d : std_logic := '0';
	
	signal bitvectord245d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled245d : std_logic := '0';
	signal matchd245d : std_logic := '0';
	
	signal bitvectord246d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled246d : std_logic := '0';
	signal matchd246d : std_logic := '0';
	
	signal bitvectord247d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled247d : std_logic := '0';
	signal matchd247d : std_logic := '0';
	
	signal bitvectord248d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled248d : std_logic := '0';
	signal matchd248d : std_logic := '0';
	
	signal bitvectord249d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled249d : std_logic := '0';
	signal matchd249d : std_logic := '0';
	
	signal bitvectord250d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled250d : std_logic := '0';
	signal matchd250d : std_logic := '0';
	
	signal bitvectord251d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled251d : std_logic := '0';
	signal matchd251d : std_logic := '0';
	
	signal bitvectord252d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled252d : std_logic := '1';
	signal matchd252d : std_logic := '0';
	
	signal bitvectord253d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled253d : std_logic := '0';
	signal matchd253d : std_logic := '0';
	
	signal bitvectord254d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled254d : std_logic := '0';
	signal matchd254d : std_logic := '0';
	
	signal bitvectord255d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled255d : std_logic := '0';
	signal matchd255d : std_logic := '0';
	
	signal bitvectord256d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled256d : std_logic := '0';
	signal matchd256d : std_logic := '0';
	
	signal bitvectord257d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled257d : std_logic := '0';
	signal matchd257d : std_logic := '0';
	
	signal bitvectord258d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled258d : std_logic := '0';
	signal matchd258d : std_logic := '0';
	
	signal bitvectord259d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled259d : std_logic := '0';
	signal matchd259d : std_logic := '0';
	
	signal bitvectord260d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled260d : std_logic := '0';
	signal matchd260d : std_logic := '0';
	
	signal bitvectord261d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled261d : std_logic := '0';
	signal matchd261d : std_logic := '0';
	
	signal bitvectord262d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled262d : std_logic := '0';
	signal matchd262d : std_logic := '0';
	
	signal bitvectord263d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled263d : std_logic := '0';
	signal matchd263d : std_logic := '0';
	
	signal bitvectord264d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled264d : std_logic := '0';
	signal matchd264d : std_logic := '0';
	
	signal bitvectord265d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled265d : std_logic := '0';
	signal matchd265d : std_logic := '0';
	
	signal bitvectord266d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled266d : std_logic := '0';
	signal matchd266d : std_logic := '0';
	
	signal bitvectord267d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled267d : std_logic := '0';
	signal matchd267d : std_logic := '0';
	
	signal bitvectord268d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled268d : std_logic := '0';
	signal matchd268d : std_logic := '0';
	
	signal bitvectord270d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled270d : std_logic := '1';
	signal matchd270d : std_logic := '0';
	
	signal bitvectord271d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled271d : std_logic := '0';
	signal matchd271d : std_logic := '0';
	
	signal bitvectord272d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled272d : std_logic := '0';
	signal matchd272d : std_logic := '0';
	
	signal bitvectord273d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled273d : std_logic := '0';
	signal matchd273d : std_logic := '0';
	
	signal bitvectord274d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled274d : std_logic := '0';
	signal matchd274d : std_logic := '0';
	
	signal bitvectord275d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled275d : std_logic := '0';
	signal matchd275d : std_logic := '0';
	
	signal bitvectord276d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled276d : std_logic := '0';
	signal matchd276d : std_logic := '0';
	
	signal bitvectord277d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled277d : std_logic := '0';
	signal matchd277d : std_logic := '0';
	
	signal bitvectord278d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled278d : std_logic := '0';
	signal matchd278d : std_logic := '0';
	
	signal bitvectord279d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled279d : std_logic := '0';
	signal matchd279d : std_logic := '0';
	
	signal bitvectord280d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled280d : std_logic := '0';
	signal matchd280d : std_logic := '0';
	
	signal bitvectord281d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled281d : std_logic := '0';
	signal matchd281d : std_logic := '0';
	
	signal bitvectord282d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled282d : std_logic := '0';
	signal matchd282d : std_logic := '0';
	
	signal bitvectord283d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled283d : std_logic := '1';
	signal matchd283d : std_logic := '0';
	
	signal bitvectord284d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled284d : std_logic := '0';
	signal matchd284d : std_logic := '0';
	
	signal bitvectord285d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled285d : std_logic := '0';
	signal matchd285d : std_logic := '0';
	
	signal bitvectord286d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled286d : std_logic := '0';
	signal matchd286d : std_logic := '0';
	
	signal bitvectord287d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled287d : std_logic := '0';
	signal matchd287d : std_logic := '0';
	
	signal bitvectord288d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled288d : std_logic := '0';
	signal matchd288d : std_logic := '0';
	
	signal bitvectord289d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled289d : std_logic := '0';
	signal matchd289d : std_logic := '0';
	
	signal bitvectord290d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled290d : std_logic := '0';
	signal matchd290d : std_logic := '0';
	
	signal bitvectord291d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled291d : std_logic := '0';
	signal matchd291d : std_logic := '0';
	
	signal bitvectord292d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled292d : std_logic := '0';
	signal matchd292d : std_logic := '0';
	
	signal bitvectord293d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled293d : std_logic := '0';
	signal matchd293d : std_logic := '0';
	
	signal bitvectord294d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled294d : std_logic := '0';
	signal matchd294d : std_logic := '0';
	
	signal bitvectord295d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled295d : std_logic := '0';
	signal matchd295d : std_logic := '0';
	
	signal bitvectord296d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled296d : std_logic := '0';
	signal matchd296d : std_logic := '0';
	
	signal bitvectord297d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled297d : std_logic := '0';
	signal matchd297d : std_logic := '0';
	
	signal bitvectord298d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled298d : std_logic := '1';
	signal matchd298d : std_logic := '0';
	
	signal bitvectord299d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled299d : std_logic := '0';
	signal matchd299d : std_logic := '0';
	
	signal bitvectord300d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled300d : std_logic := '0';
	signal matchd300d : std_logic := '0';
	
	signal bitvectord301d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled301d : std_logic := '0';
	signal matchd301d : std_logic := '0';
	
	signal bitvectord302d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled302d : std_logic := '0';
	signal matchd302d : std_logic := '0';
	
	signal bitvectord303d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled303d : std_logic := '0';
	signal matchd303d : std_logic := '0';
	
	signal bitvectord304d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled304d : std_logic := '0';
	signal matchd304d : std_logic := '0';
	
	signal bitvectord305d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled305d : std_logic := '0';
	signal matchd305d : std_logic := '0';
	
	signal bitvectord306d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled306d : std_logic := '0';
	signal matchd306d : std_logic := '0';
	
	signal bitvectord307d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled307d : std_logic := '0';
	signal matchd307d : std_logic := '0';
	
	signal bitvectord308d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled308d : std_logic := '0';
	signal matchd308d : std_logic := '0';
	
	signal bitvectord309d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled309d : std_logic := '0';
	signal matchd309d : std_logic := '0';
	
	signal bitvectord310d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled310d : std_logic := '0';
	signal matchd310d : std_logic := '0';
	
	signal bitvectord311d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled311d : std_logic := '0';
	signal matchd311d : std_logic := '0';
	
	signal bitvectord312d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled312d : std_logic := '0';
	signal matchd312d : std_logic := '0';
	
	signal bitvectord314d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled314d : std_logic := '1';
	signal matchd314d : std_logic := '0';
	
	signal bitvectord315d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled315d : std_logic := '0';
	signal matchd315d : std_logic := '0';
	
	signal bitvectord316d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled316d : std_logic := '0';
	signal matchd316d : std_logic := '0';
	
	signal bitvectord317d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled317d : std_logic := '0';
	signal matchd317d : std_logic := '0';
	
	signal bitvectord318d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled318d : std_logic := '0';
	signal matchd318d : std_logic := '0';
	
	signal bitvectord319d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled319d : std_logic := '0';
	signal matchd319d : std_logic := '0';
	
	signal bitvectord320d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled320d : std_logic := '0';
	signal matchd320d : std_logic := '0';
	
	signal bitvectord321d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled321d : std_logic := '0';
	signal matchd321d : std_logic := '0';
	
	signal bitvectord322d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled322d : std_logic := '0';
	signal matchd322d : std_logic := '0';
	
	signal bitvectord323d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled323d : std_logic := '0';
	signal matchd323d : std_logic := '0';
	
	signal bitvectord324d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled324d : std_logic := '0';
	signal matchd324d : std_logic := '0';
	
	signal bitvectord325d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled325d : std_logic := '0';
	signal matchd325d : std_logic := '0';
	
	signal bitvectord326d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled326d : std_logic := '1';
	signal matchd326d : std_logic := '0';
	
	signal bitvectord327d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled327d : std_logic := '0';
	signal matchd327d : std_logic := '0';
	
	signal bitvectord328d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled328d : std_logic := '0';
	signal matchd328d : std_logic := '0';
	
	signal bitvectord329d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled329d : std_logic := '0';
	signal matchd329d : std_logic := '0';
	
	signal bitvectord330d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled330d : std_logic := '0';
	signal matchd330d : std_logic := '0';
	
	signal bitvectord331d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled331d : std_logic := '0';
	signal matchd331d : std_logic := '0';
	
	signal bitvectord332d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled332d : std_logic := '0';
	signal matchd332d : std_logic := '0';
	
	signal bitvectord333d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled333d : std_logic := '0';
	signal matchd333d : std_logic := '0';
	
	signal bitvectord334d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled334d : std_logic := '0';
	signal matchd334d : std_logic := '0';
	
	signal bitvectord335d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled335d : std_logic := '0';
	signal matchd335d : std_logic := '0';
	
	signal bitvectord336d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled336d : std_logic := '0';
	signal matchd336d : std_logic := '0';
	
	signal bitvectord337d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled337d : std_logic := '0';
	signal matchd337d : std_logic := '0';
	
	signal bitvectord338d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled338d : std_logic := '0';
	signal matchd338d : std_logic := '0';
	
	signal bitvectord339d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled339d : std_logic := '0';
	signal matchd339d : std_logic := '0';
	
	signal bitvectord340d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled340d : std_logic := '0';
	signal matchd340d : std_logic := '0';
	
	signal bitvectord341d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled341d : std_logic := '1';
	signal matchd341d : std_logic := '0';
	
	signal bitvectord342d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled342d : std_logic := '0';
	signal matchd342d : std_logic := '0';
	
	signal bitvectord343d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled343d : std_logic := '0';
	signal matchd343d : std_logic := '0';
	
	signal bitvectord344d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled344d : std_logic := '0';
	signal matchd344d : std_logic := '0';
	
	signal bitvectord345d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled345d : std_logic := '0';
	signal matchd345d : std_logic := '0';
	
	signal bitvectord346d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled346d : std_logic := '0';
	signal matchd346d : std_logic := '0';
	
	signal bitvectord347d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled347d : std_logic := '0';
	signal matchd347d : std_logic := '0';
	
	signal bitvectord348d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled348d : std_logic := '0';
	signal matchd348d : std_logic := '0';
	
	signal bitvectord349d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled349d : std_logic := '0';
	signal matchd349d : std_logic := '0';
	
	signal bitvectord350d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled350d : std_logic := '0';
	signal matchd350d : std_logic := '0';
	
	signal bitvectord351d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled351d : std_logic := '0';
	signal matchd351d : std_logic := '0';
	
	signal bitvectord352d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled352d : std_logic := '0';
	signal matchd352d : std_logic := '0';
	
	signal bitvectord353d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled353d : std_logic := '0';
	signal matchd353d : std_logic := '0';
	
	signal bitvectord354d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled354d : std_logic := '0';
	signal matchd354d : std_logic := '0';
	
	signal bitvectord355d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled355d : std_logic := '0';
	signal matchd355d : std_logic := '0';
	
	signal bitvectord357d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled357d : std_logic := '1';
	signal matchd357d : std_logic := '0';
	
	signal bitvectord358d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled358d : std_logic := '0';
	signal matchd358d : std_logic := '0';
	
	signal bitvectord359d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled359d : std_logic := '0';
	signal matchd359d : std_logic := '0';
	
	signal bitvectord360d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled360d : std_logic := '0';
	signal matchd360d : std_logic := '0';
	
	signal bitvectord361d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled361d : std_logic := '0';
	signal matchd361d : std_logic := '0';
	
	signal bitvectord362d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled362d : std_logic := '0';
	signal matchd362d : std_logic := '0';
	
	signal bitvectord363d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled363d : std_logic := '0';
	signal matchd363d : std_logic := '0';
	
	signal bitvectord364d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled364d : std_logic := '0';
	signal matchd364d : std_logic := '0';
	
	signal bitvectord365d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled365d : std_logic := '0';
	signal matchd365d : std_logic := '0';
	
	signal bitvectord366d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled366d : std_logic := '0';
	signal matchd366d : std_logic := '0';
	
	signal bitvectord367d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled367d : std_logic := '0';
	signal matchd367d : std_logic := '0';
	
	signal bitvectord368d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled368d : std_logic := '0';
	signal matchd368d : std_logic := '0';
	
	signal bitvectord369d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled369d : std_logic := '0';
	signal matchd369d : std_logic := '0';
	
	signal bitvectord370d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled370d : std_logic := '1';
	signal matchd370d : std_logic := '0';
	
	signal bitvectord371d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled371d : std_logic := '0';
	signal matchd371d : std_logic := '0';
	
	signal bitvectord372d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled372d : std_logic := '0';
	signal matchd372d : std_logic := '0';
	
	signal bitvectord373d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled373d : std_logic := '0';
	signal matchd373d : std_logic := '0';
	
	signal bitvectord374d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled374d : std_logic := '0';
	signal matchd374d : std_logic := '0';
	
	signal bitvectord375d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled375d : std_logic := '0';
	signal matchd375d : std_logic := '0';
	
	signal bitvectord376d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled376d : std_logic := '0';
	signal matchd376d : std_logic := '0';
	
	signal bitvectord377d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled377d : std_logic := '0';
	signal matchd377d : std_logic := '0';
	
	signal bitvectord378d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled378d : std_logic := '0';
	signal matchd378d : std_logic := '0';
	
	signal bitvectord379d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled379d : std_logic := '0';
	signal matchd379d : std_logic := '0';
	
	signal bitvectord380d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled380d : std_logic := '0';
	signal matchd380d : std_logic := '0';
	
	signal bitvectord381d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled381d : std_logic := '0';
	signal matchd381d : std_logic := '0';
	
	signal bitvectord382d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled382d : std_logic := '0';
	signal matchd382d : std_logic := '0';
	
	signal bitvectord383d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled383d : std_logic := '0';
	signal matchd383d : std_logic := '0';
	
	signal bitvectord384d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled384d : std_logic := '0';
	signal matchd384d : std_logic := '0';
	
	signal bitvectord385d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled385d : std_logic := '0';
	signal matchd385d : std_logic := '0';
	
	signal bitvectord386d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled386d : std_logic := '0';
	signal matchd386d : std_logic := '0';
	
	signal bitvectord387d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled387d : std_logic := '0';
	signal matchd387d : std_logic := '0';
	
	signal bitvectord388d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled388d : std_logic := '0';
	signal matchd388d : std_logic := '0';
	
	signal bitvectord389d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled389d : std_logic := '0';
	signal matchd389d : std_logic := '0';
	
	signal bitvectord390d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled390d : std_logic := '0';
	signal matchd390d : std_logic := '0';
	
	signal bitvectord391d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled391d : std_logic := '1';
	signal matchd391d : std_logic := '0';
	
	signal bitvectord392d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled392d : std_logic := '0';
	signal matchd392d : std_logic := '0';
	
	signal bitvectord393d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled393d : std_logic := '0';
	signal matchd393d : std_logic := '0';
	
	signal bitvectord394d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled394d : std_logic := '0';
	signal matchd394d : std_logic := '0';
	
	signal bitvectord395d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled395d : std_logic := '0';
	signal matchd395d : std_logic := '0';
	
	signal bitvectord396d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled396d : std_logic := '0';
	signal matchd396d : std_logic := '0';
	
	signal bitvectord397d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled397d : std_logic := '0';
	signal matchd397d : std_logic := '0';
	
	signal bitvectord398d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled398d : std_logic := '0';
	signal matchd398d : std_logic := '0';
	
	signal bitvectord399d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled399d : std_logic := '0';
	signal matchd399d : std_logic := '0';
	
	signal bitvectord400d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled400d : std_logic := '0';
	signal matchd400d : std_logic := '0';
	
	signal bitvectord401d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled401d : std_logic := '0';
	signal matchd401d : std_logic := '0';
	
	signal bitvectord402d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled402d : std_logic := '0';
	signal matchd402d : std_logic := '0';
	
	signal bitvectord403d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled403d : std_logic := '0';
	signal matchd403d : std_logic := '0';
	
	signal bitvectord404d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled404d : std_logic := '0';
	signal matchd404d : std_logic := '0';
	
	signal bitvectord405d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled405d : std_logic := '0';
	signal matchd405d : std_logic := '0';
	
	signal bitvectord406d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled406d : std_logic := '0';
	signal matchd406d : std_logic := '0';
	
	signal bitvectord407d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled407d : std_logic := '0';
	signal matchd407d : std_logic := '0';
	
	signal bitvectord408d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled408d : std_logic := '0';
	signal matchd408d : std_logic := '0';
	
	signal bitvectord409d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled409d : std_logic := '0';
	signal matchd409d : std_logic := '0';
	
	signal bitvectord410d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled410d : std_logic := '0';
	signal matchd410d : std_logic := '0';
	
	signal bitvectord411d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled411d : std_logic := '0';
	signal matchd411d : std_logic := '0';
	
	signal bitvectord412d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled412d : std_logic := '1';
	signal matchd412d : std_logic := '0';
	
	signal bitvectord413d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled413d : std_logic := '0';
	signal matchd413d : std_logic := '0';
	
	signal bitvectord414d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled414d : std_logic := '0';
	signal matchd414d : std_logic := '0';
	
	signal bitvectord415d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled415d : std_logic := '0';
	signal matchd415d : std_logic := '0';
	
	signal bitvectord416d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled416d : std_logic := '0';
	signal matchd416d : std_logic := '0';
	
	signal bitvectord417d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled417d : std_logic := '0';
	signal matchd417d : std_logic := '0';
	
	signal bitvectord418d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled418d : std_logic := '0';
	signal matchd418d : std_logic := '0';
	
	signal bitvectord419d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled419d : std_logic := '0';
	signal matchd419d : std_logic := '0';
	
	signal bitvectord420d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled420d : std_logic := '0';
	signal matchd420d : std_logic := '0';
	
	signal bitvectord421d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled421d : std_logic := '0';
	signal matchd421d : std_logic := '0';
	
	signal bitvectord422d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled422d : std_logic := '0';
	signal matchd422d : std_logic := '0';
	
	signal bitvectord423d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled423d : std_logic := '0';
	signal matchd423d : std_logic := '0';
	
	signal bitvectord424d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled424d : std_logic := '0';
	signal matchd424d : std_logic := '0';
	
	signal bitvectord425d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled425d : std_logic := '0';
	signal matchd425d : std_logic := '0';
	
	signal bitvectord426d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled426d : std_logic := '0';
	signal matchd426d : std_logic := '0';
	
	signal bitvectord427d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled427d : std_logic := '0';
	signal matchd427d : std_logic := '0';
	
	signal bitvectord428d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled428d : std_logic := '0';
	signal matchd428d : std_logic := '0';
	
	signal bitvectord429d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled429d : std_logic := '0';
	signal matchd429d : std_logic := '0';
	
	signal bitvectord430d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled430d : std_logic := '0';
	signal matchd430d : std_logic := '0';
	
	signal bitvectord431d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled431d : std_logic := '0';
	signal matchd431d : std_logic := '0';
	
	signal bitvectord432d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled432d : std_logic := '0';
	signal matchd432d : std_logic := '0';
	
	signal bitvectord434d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled434d : std_logic := '1';
	signal matchd434d : std_logic := '0';
	
	signal bitvectord435d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled435d : std_logic := '0';
	signal matchd435d : std_logic := '0';
	
	signal bitvectord436d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled436d : std_logic := '0';
	signal matchd436d : std_logic := '0';
	
	signal bitvectord437d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled437d : std_logic := '0';
	signal matchd437d : std_logic := '0';
	
	signal bitvectord438d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled438d : std_logic := '0';
	signal matchd438d : std_logic := '0';
	
	signal bitvectord439d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled439d : std_logic := '0';
	signal matchd439d : std_logic := '0';
	
	signal bitvectord440d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled440d : std_logic := '0';
	signal matchd440d : std_logic := '0';
	
	signal bitvectord441d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled441d : std_logic := '0';
	signal matchd441d : std_logic := '0';
	
	signal bitvectord442d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled442d : std_logic := '0';
	signal matchd442d : std_logic := '0';
	
	signal bitvectord443d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled443d : std_logic := '0';
	signal matchd443d : std_logic := '0';
	
	signal bitvectord444d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled444d : std_logic := '0';
	signal matchd444d : std_logic := '0';
	
	signal bitvectord445d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled445d : std_logic := '1';
	signal matchd445d : std_logic := '0';
	
	signal bitvectord446d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled446d : std_logic := '0';
	signal matchd446d : std_logic := '0';
	
	signal bitvectord447d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled447d : std_logic := '0';
	signal matchd447d : std_logic := '0';
	
	signal bitvectord448d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled448d : std_logic := '0';
	signal matchd448d : std_logic := '0';
	
	signal bitvectord449d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled449d : std_logic := '0';
	signal matchd449d : std_logic := '0';
	
	signal bitvectord450d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled450d : std_logic := '0';
	signal matchd450d : std_logic := '0';
	
	signal bitvectord451d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled451d : std_logic := '0';
	signal matchd451d : std_logic := '0';
	
	signal bitvectord452d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled452d : std_logic := '0';
	signal matchd452d : std_logic := '0';
	
	signal bitvectord453d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled453d : std_logic := '0';
	signal matchd453d : std_logic := '0';
	
	signal bitvectord454d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled454d : std_logic := '0';
	signal matchd454d : std_logic := '0';
	
	signal bitvectord455d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled455d : std_logic := '0';
	signal matchd455d : std_logic := '0';
	
	signal bitvectord456d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled456d : std_logic := '0';
	signal matchd456d : std_logic := '0';
	
	signal bitvectord457d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled457d : std_logic := '0';
	signal matchd457d : std_logic := '0';
	
	signal bitvectord458d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled458d : std_logic := '0';
	signal matchd458d : std_logic := '0';
	
	signal bitvectord459d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled459d : std_logic := '0';
	signal matchd459d : std_logic := '0';
	
	signal bitvectord460d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled460d : std_logic := '0';
	signal matchd460d : std_logic := '0';
	
	signal bitvectord461d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled461d : std_logic := '0';
	signal matchd461d : std_logic := '0';
	
	signal bitvectord462d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled462d : std_logic := '0';
	signal matchd462d : std_logic := '0';
	
	signal bitvectord463d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled463d : std_logic := '0';
	signal matchd463d : std_logic := '0';
	
	signal bitvectord464d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled464d : std_logic := '0';
	signal matchd464d : std_logic := '0';
	
	signal bitvectord465d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled465d : std_logic := '1';
	signal matchd465d : std_logic := '0';
	
	signal bitvectord466d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled466d : std_logic := '0';
	signal matchd466d : std_logic := '0';
	
	signal bitvectord467d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled467d : std_logic := '0';
	signal matchd467d : std_logic := '0';
	
	signal bitvectord468d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled468d : std_logic := '0';
	signal matchd468d : std_logic := '0';
	
	signal bitvectord469d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled469d : std_logic := '0';
	signal matchd469d : std_logic := '0';
	
	signal bitvectord470d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled470d : std_logic := '0';
	signal matchd470d : std_logic := '0';
	
	signal bitvectord471d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled471d : std_logic := '0';
	signal matchd471d : std_logic := '0';
	
	signal bitvectord472d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled472d : std_logic := '0';
	signal matchd472d : std_logic := '0';
	
	signal bitvectord473d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled473d : std_logic := '0';
	signal matchd473d : std_logic := '0';
	
	signal bitvectord474d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled474d : std_logic := '0';
	signal matchd474d : std_logic := '0';
	
	signal bitvectord475d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled475d : std_logic := '0';
	signal matchd475d : std_logic := '0';
	
	signal bitvectord476d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled476d : std_logic := '0';
	signal matchd476d : std_logic := '0';
	
	signal bitvectord477d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled477d : std_logic := '0';
	signal matchd477d : std_logic := '0';
	
	signal bitvectord478d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled478d : std_logic := '0';
	signal matchd478d : std_logic := '0';
	
	signal bitvectord479d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled479d : std_logic := '0';
	signal matchd479d : std_logic := '0';
	
	signal bitvectord480d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled480d : std_logic := '0';
	signal matchd480d : std_logic := '0';
	
	signal bitvectord481d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled481d : std_logic := '0';
	signal matchd481d : std_logic := '0';
	
	signal bitvectord482d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled482d : std_logic := '0';
	signal matchd482d : std_logic := '0';
	
	signal bitvectord483d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled483d : std_logic := '0';
	signal matchd483d : std_logic := '0';
	
	signal bitvectord484d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled484d : std_logic := '0';
	signal matchd484d : std_logic := '0';
	
	signal bitvectord485d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled485d : std_logic := '1';
	signal matchd485d : std_logic := '0';
	
	signal bitvectord486d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled486d : std_logic := '0';
	signal matchd486d : std_logic := '0';
	
	signal bitvectord487d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled487d : std_logic := '0';
	signal matchd487d : std_logic := '0';
	
	signal bitvectord488d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled488d : std_logic := '0';
	signal matchd488d : std_logic := '0';
	
	signal bitvectord489d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled489d : std_logic := '0';
	signal matchd489d : std_logic := '0';
	
	signal bitvectord490d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled490d : std_logic := '0';
	signal matchd490d : std_logic := '0';
	
	signal bitvectord491d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled491d : std_logic := '0';
	signal matchd491d : std_logic := '0';
	
	signal bitvectord492d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled492d : std_logic := '0';
	signal matchd492d : std_logic := '0';
	
	signal bitvectord493d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled493d : std_logic := '0';
	signal matchd493d : std_logic := '0';
	
	signal bitvectord494d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled494d : std_logic := '0';
	signal matchd494d : std_logic := '0';
	
	signal bitvectord495d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled495d : std_logic := '0';
	signal matchd495d : std_logic := '0';
	
	signal bitvectord496d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled496d : std_logic := '0';
	signal matchd496d : std_logic := '0';
	
	signal bitvectord497d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled497d : std_logic := '0';
	signal matchd497d : std_logic := '0';
	
	signal bitvectord498d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled498d : std_logic := '0';
	signal matchd498d : std_logic := '0';
	
	signal bitvectord499d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled499d : std_logic := '0';
	signal matchd499d : std_logic := '0';
	
	signal bitvectord500d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled500d : std_logic := '0';
	signal matchd500d : std_logic := '0';
	
	signal bitvectord501d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled501d : std_logic := '0';
	signal matchd501d : std_logic := '0';
	
	signal bitvectord502d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled502d : std_logic := '0';
	signal matchd502d : std_logic := '0';
	
	signal bitvectord503d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled503d : std_logic := '0';
	signal matchd503d : std_logic := '0';
	
	signal bitvectord504d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled504d : std_logic := '0';
	signal matchd504d : std_logic := '0';
	
	signal bitvectord506d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled506d : std_logic := '1';
	signal matchd506d : std_logic := '0';
	
	signal bitvectord507d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled507d : std_logic := '0';
	signal matchd507d : std_logic := '0';
	
	signal bitvectord508d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled508d : std_logic := '0';
	signal matchd508d : std_logic := '0';
	
	signal bitvectord509d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled509d : std_logic := '0';
	signal matchd509d : std_logic := '0';
	
	signal bitvectord510d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled510d : std_logic := '0';
	signal matchd510d : std_logic := '0';
	
	signal bitvectord511d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled511d : std_logic := '0';
	signal matchd511d : std_logic := '0';
	
	signal bitvectord512d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled512d : std_logic := '0';
	signal matchd512d : std_logic := '0';
	
	signal bitvectord513d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled513d : std_logic := '0';
	signal matchd513d : std_logic := '0';
	
	signal bitvectord514d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled514d : std_logic := '0';
	signal matchd514d : std_logic := '0';
	
	signal bitvectord515d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled515d : std_logic := '0';
	signal matchd515d : std_logic := '0';
	
	signal bitvectord516d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled516d : std_logic := '0';
	signal matchd516d : std_logic := '0';
	
	signal bitvectord517d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled517d : std_logic := '0';
	signal matchd517d : std_logic := '0';
	
	signal bitvectord518d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled518d : std_logic := '0';
	signal matchd518d : std_logic := '0';
	
	signal bitvectord519d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled519d : std_logic := '0';
	signal matchd519d : std_logic := '0';
	
	signal bitvectord520d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled520d : std_logic := '0';
	signal matchd520d : std_logic := '0';
	
	signal bitvectord521d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled521d : std_logic := '0';
	signal matchd521d : std_logic := '0';
	
	signal bitvectord522d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled522d : std_logic := '1';
	signal matchd522d : std_logic := '0';
	
	signal bitvectord523d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled523d : std_logic := '0';
	signal matchd523d : std_logic := '0';
	
	signal bitvectord524d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled524d : std_logic := '0';
	signal matchd524d : std_logic := '0';
	
	signal bitvectord525d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled525d : std_logic := '0';
	signal matchd525d : std_logic := '0';
	
	signal bitvectord526d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled526d : std_logic := '0';
	signal matchd526d : std_logic := '0';
	
	signal bitvectord527d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled527d : std_logic := '0';
	signal matchd527d : std_logic := '0';
	
	signal bitvectord528d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled528d : std_logic := '0';
	signal matchd528d : std_logic := '0';
	
	signal bitvectord529d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled529d : std_logic := '0';
	signal matchd529d : std_logic := '0';
	
	signal bitvectord530d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled530d : std_logic := '0';
	signal matchd530d : std_logic := '0';
	
	signal bitvectord531d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled531d : std_logic := '0';
	signal matchd531d : std_logic := '0';
	
	signal bitvectord532d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled532d : std_logic := '0';
	signal matchd532d : std_logic := '0';
	
	signal bitvectord533d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled533d : std_logic := '0';
	signal matchd533d : std_logic := '0';
	
	signal bitvectord534d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled534d : std_logic := '0';
	signal matchd534d : std_logic := '0';
	
	signal bitvectord535d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled535d : std_logic := '0';
	signal matchd535d : std_logic := '0';
	
	signal bitvectord536d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled536d : std_logic := '0';
	signal matchd536d : std_logic := '0';
	
	signal bitvectord537d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled537d : std_logic := '0';
	signal matchd537d : std_logic := '0';
	
	signal bitvectord538d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled538d : std_logic := '1';
	signal matchd538d : std_logic := '0';
	
	signal bitvectord539d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled539d : std_logic := '0';
	signal matchd539d : std_logic := '0';
	
	signal bitvectord540d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled540d : std_logic := '0';
	signal matchd540d : std_logic := '0';
	
	signal bitvectord541d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled541d : std_logic := '0';
	signal matchd541d : std_logic := '0';
	
	signal bitvectord542d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled542d : std_logic := '0';
	signal matchd542d : std_logic := '0';
	
	signal bitvectord543d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled543d : std_logic := '0';
	signal matchd543d : std_logic := '0';
	
	signal bitvectord544d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled544d : std_logic := '0';
	signal matchd544d : std_logic := '0';
	
	signal bitvectord545d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled545d : std_logic := '0';
	signal matchd545d : std_logic := '0';
	
	signal bitvectord546d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled546d : std_logic := '0';
	signal matchd546d : std_logic := '0';
	
	signal bitvectord547d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled547d : std_logic := '0';
	signal matchd547d : std_logic := '0';
	
	signal bitvectord548d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled548d : std_logic := '0';
	signal matchd548d : std_logic := '0';
	
	signal bitvectord549d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled549d : std_logic := '0';
	signal matchd549d : std_logic := '0';
	
	signal bitvectord550d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled550d : std_logic := '0';
	signal matchd550d : std_logic := '0';
	
	signal bitvectord551d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled551d : std_logic := '0';
	signal matchd551d : std_logic := '0';
	
	signal bitvectord552d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled552d : std_logic := '0';
	signal matchd552d : std_logic := '0';
	
	signal bitvectord553d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled553d : std_logic := '0';
	signal matchd553d : std_logic := '0';
	
	signal bitvectord555d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled555d : std_logic := '1';
	signal matchd555d : std_logic := '0';
	
	signal bitvectord556d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled556d : std_logic := '0';
	signal matchd556d : std_logic := '0';
	
	signal bitvectord557d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled557d : std_logic := '0';
	signal matchd557d : std_logic := '0';
	
	signal bitvectord558d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled558d : std_logic := '0';
	signal matchd558d : std_logic := '0';
	
	signal bitvectord559d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled559d : std_logic := '0';
	signal matchd559d : std_logic := '0';
	
	signal bitvectord560d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled560d : std_logic := '0';
	signal matchd560d : std_logic := '0';
	
	signal bitvectord561d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled561d : std_logic := '0';
	signal matchd561d : std_logic := '0';
	
	signal bitvectord562d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled562d : std_logic := '0';
	signal matchd562d : std_logic := '0';
	
	signal bitvectord563d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled563d : std_logic := '0';
	signal matchd563d : std_logic := '0';
	
	signal bitvectord564d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled564d : std_logic := '0';
	signal matchd564d : std_logic := '0';
	
	signal bitvectord565d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled565d : std_logic := '0';
	signal matchd565d : std_logic := '0';
	
	signal bitvectord566d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled566d : std_logic := '1';
	signal matchd566d : std_logic := '0';
	
	signal bitvectord567d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled567d : std_logic := '0';
	signal matchd567d : std_logic := '0';
	
	signal bitvectord568d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled568d : std_logic := '0';
	signal matchd568d : std_logic := '0';
	
	signal bitvectord569d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled569d : std_logic := '0';
	signal matchd569d : std_logic := '0';
	
	signal bitvectord570d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled570d : std_logic := '0';
	signal matchd570d : std_logic := '0';
	
	signal bitvectord571d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled571d : std_logic := '0';
	signal matchd571d : std_logic := '0';
	
	signal bitvectord572d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled572d : std_logic := '0';
	signal matchd572d : std_logic := '0';
	
	signal bitvectord573d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled573d : std_logic := '0';
	signal matchd573d : std_logic := '0';
	
	signal bitvectord574d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled574d : std_logic := '0';
	signal matchd574d : std_logic := '0';
	
	signal bitvectord575d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled575d : std_logic := '0';
	signal matchd575d : std_logic := '0';
	
	signal bitvectord576d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled576d : std_logic := '0';
	signal matchd576d : std_logic := '0';
	
	signal bitvectord577d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled577d : std_logic := '0';
	signal matchd577d : std_logic := '0';
	
	signal bitvectord578d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled578d : std_logic := '0';
	signal matchd578d : std_logic := '0';
	
	signal bitvectord579d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled579d : std_logic := '0';
	signal matchd579d : std_logic := '0';
	
	signal bitvectord580d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled580d : std_logic := '0';
	signal matchd580d : std_logic := '0';
	
	signal bitvectord581d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled581d : std_logic := '0';
	signal matchd581d : std_logic := '0';
	
	signal bitvectord582d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled582d : std_logic := '0';
	signal matchd582d : std_logic := '0';
	
	signal bitvectord583d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled583d : std_logic := '0';
	signal matchd583d : std_logic := '0';
	
	signal bitvectord584d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled584d : std_logic := '0';
	signal matchd584d : std_logic := '0';
	
	signal bitvectord585d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled585d : std_logic := '0';
	signal matchd585d : std_logic := '0';
	
	signal bitvectord586d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled586d : std_logic := '1';
	signal matchd586d : std_logic := '0';
	
	signal bitvectord587d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled587d : std_logic := '0';
	signal matchd587d : std_logic := '0';
	
	signal bitvectord588d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled588d : std_logic := '0';
	signal matchd588d : std_logic := '0';
	
	signal bitvectord589d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled589d : std_logic := '0';
	signal matchd589d : std_logic := '0';
	
	signal bitvectord590d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled590d : std_logic := '0';
	signal matchd590d : std_logic := '0';
	
	signal bitvectord591d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled591d : std_logic := '0';
	signal matchd591d : std_logic := '0';
	
	signal bitvectord592d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled592d : std_logic := '0';
	signal matchd592d : std_logic := '0';
	
	signal bitvectord593d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled593d : std_logic := '0';
	signal matchd593d : std_logic := '0';
	
	signal bitvectord594d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled594d : std_logic := '0';
	signal matchd594d : std_logic := '0';
	
	signal bitvectord595d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled595d : std_logic := '0';
	signal matchd595d : std_logic := '0';
	
	signal bitvectord596d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled596d : std_logic := '0';
	signal matchd596d : std_logic := '0';
	
	signal bitvectord597d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled597d : std_logic := '0';
	signal matchd597d : std_logic := '0';
	
	signal bitvectord598d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled598d : std_logic := '0';
	signal matchd598d : std_logic := '0';
	
	signal bitvectord599d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled599d : std_logic := '0';
	signal matchd599d : std_logic := '0';
	
	signal bitvectord600d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled600d : std_logic := '0';
	signal matchd600d : std_logic := '0';
	
	signal bitvectord601d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled601d : std_logic := '0';
	signal matchd601d : std_logic := '0';
	
	signal bitvectord602d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled602d : std_logic := '0';
	signal matchd602d : std_logic := '0';
	
	signal bitvectord603d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled603d : std_logic := '0';
	signal matchd603d : std_logic := '0';
	
	signal bitvectord604d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled604d : std_logic := '0';
	signal matchd604d : std_logic := '0';
	
	signal bitvectord605d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled605d : std_logic := '0';
	signal matchd605d : std_logic := '0';
	
	signal bitvectord606d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled606d : std_logic := '1';
	signal matchd606d : std_logic := '0';
	
	signal bitvectord607d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled607d : std_logic := '0';
	signal matchd607d : std_logic := '0';
	
	signal bitvectord608d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled608d : std_logic := '0';
	signal matchd608d : std_logic := '0';
	
	signal bitvectord609d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled609d : std_logic := '0';
	signal matchd609d : std_logic := '0';
	
	signal bitvectord610d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled610d : std_logic := '0';
	signal matchd610d : std_logic := '0';
	
	signal bitvectord611d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled611d : std_logic := '0';
	signal matchd611d : std_logic := '0';
	
	signal bitvectord612d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled612d : std_logic := '0';
	signal matchd612d : std_logic := '0';
	
	signal bitvectord613d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled613d : std_logic := '0';
	signal matchd613d : std_logic := '0';
	
	signal bitvectord614d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled614d : std_logic := '0';
	signal matchd614d : std_logic := '0';
	
	signal bitvectord615d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled615d : std_logic := '0';
	signal matchd615d : std_logic := '0';
	
	signal bitvectord616d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled616d : std_logic := '0';
	signal matchd616d : std_logic := '0';
	
	signal bitvectord617d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled617d : std_logic := '0';
	signal matchd617d : std_logic := '0';
	
	signal bitvectord618d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled618d : std_logic := '0';
	signal matchd618d : std_logic := '0';
	
	signal bitvectord619d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled619d : std_logic := '0';
	signal matchd619d : std_logic := '0';
	
	signal bitvectord620d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled620d : std_logic := '0';
	signal matchd620d : std_logic := '0';
	
	signal bitvectord621d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled621d : std_logic := '0';
	signal matchd621d : std_logic := '0';
	
	signal bitvectord622d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled622d : std_logic := '0';
	signal matchd622d : std_logic := '0';
	
	signal bitvectord623d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled623d : std_logic := '0';
	signal matchd623d : std_logic := '0';
	
	signal bitvectord624d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled624d : std_logic := '0';
	signal matchd624d : std_logic := '0';
	
	signal bitvectord625d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled625d : std_logic := '0';
	signal matchd625d : std_logic := '0';
	
	signal bitvectord627d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled627d : std_logic := '1';
	signal matchd627d : std_logic := '0';
	
	signal bitvectord628d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled628d : std_logic := '0';
	signal matchd628d : std_logic := '0';
	
	signal bitvectord629d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled629d : std_logic := '0';
	signal matchd629d : std_logic := '0';
	
	signal bitvectord630d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled630d : std_logic := '0';
	signal matchd630d : std_logic := '0';
	
	signal bitvectord631d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled631d : std_logic := '0';
	signal matchd631d : std_logic := '0';
	
	signal bitvectord632d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled632d : std_logic := '0';
	signal matchd632d : std_logic := '0';
	
	signal bitvectord633d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled633d : std_logic := '0';
	signal matchd633d : std_logic := '0';
	
	signal bitvectord634d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled634d : std_logic := '0';
	signal matchd634d : std_logic := '0';
	
	signal bitvectord635d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled635d : std_logic := '0';
	signal matchd635d : std_logic := '0';
	
	signal bitvectord636d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled636d : std_logic := '0';
	signal matchd636d : std_logic := '0';
	
	signal bitvectord637d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled637d : std_logic := '0';
	signal matchd637d : std_logic := '0';
	
	signal bitvectord638d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled638d : std_logic := '0';
	signal matchd638d : std_logic := '0';
	
	signal bitvectord639d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled639d : std_logic := '0';
	signal matchd639d : std_logic := '0';
	
	signal bitvectord640d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled640d : std_logic := '1';
	signal matchd640d : std_logic := '0';
	
	signal bitvectord641d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled641d : std_logic := '0';
	signal matchd641d : std_logic := '0';
	
	signal bitvectord642d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled642d : std_logic := '0';
	signal matchd642d : std_logic := '0';
	
	signal bitvectord643d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled643d : std_logic := '0';
	signal matchd643d : std_logic := '0';
	
	signal bitvectord644d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled644d : std_logic := '0';
	signal matchd644d : std_logic := '0';
	
	signal bitvectord645d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled645d : std_logic := '0';
	signal matchd645d : std_logic := '0';
	
	signal bitvectord646d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled646d : std_logic := '0';
	signal matchd646d : std_logic := '0';
	
	signal bitvectord647d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled647d : std_logic := '0';
	signal matchd647d : std_logic := '0';
	
	signal bitvectord648d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled648d : std_logic := '0';
	signal matchd648d : std_logic := '0';
	
	signal bitvectord649d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled649d : std_logic := '0';
	signal matchd649d : std_logic := '0';
	
	signal bitvectord650d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled650d : std_logic := '0';
	signal matchd650d : std_logic := '0';
	
	signal bitvectord651d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled651d : std_logic := '0';
	signal matchd651d : std_logic := '0';
	
	signal bitvectord652d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled652d : std_logic := '1';
	signal matchd652d : std_logic := '0';
	
	signal bitvectord653d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled653d : std_logic := '0';
	signal matchd653d : std_logic := '0';
	
	signal bitvectord654d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled654d : std_logic := '0';
	signal matchd654d : std_logic := '0';
	
	signal bitvectord655d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled655d : std_logic := '0';
	signal matchd655d : std_logic := '0';
	
	signal bitvectord656d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled656d : std_logic := '0';
	signal matchd656d : std_logic := '0';
	
	signal bitvectord657d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled657d : std_logic := '0';
	signal matchd657d : std_logic := '0';
	
	signal bitvectord658d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled658d : std_logic := '0';
	signal matchd658d : std_logic := '0';
	
	signal bitvectord659d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled659d : std_logic := '0';
	signal matchd659d : std_logic := '0';
	
	signal bitvectord660d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled660d : std_logic := '0';
	signal matchd660d : std_logic := '0';
	
	signal bitvectord661d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled661d : std_logic := '0';
	signal matchd661d : std_logic := '0';
	
	signal bitvectord662d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled662d : std_logic := '0';
	signal matchd662d : std_logic := '0';
	
	signal bitvectord663d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled663d : std_logic := '1';
	signal matchd663d : std_logic := '0';
	
	signal bitvectord664d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled664d : std_logic := '0';
	signal matchd664d : std_logic := '0';
	
	signal bitvectord665d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled665d : std_logic := '0';
	signal matchd665d : std_logic := '0';
	
	signal bitvectord666d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled666d : std_logic := '0';
	signal matchd666d : std_logic := '0';
	
	signal bitvectord667d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled667d : std_logic := '0';
	signal matchd667d : std_logic := '0';
	
	signal bitvectord668d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled668d : std_logic := '0';
	signal matchd668d : std_logic := '0';
	
	signal bitvectord669d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled669d : std_logic := '0';
	signal matchd669d : std_logic := '0';
	
	signal bitvectord670d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled670d : std_logic := '0';
	signal matchd670d : std_logic := '0';
	
	signal bitvectord671d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled671d : std_logic := '0';
	signal matchd671d : std_logic := '0';
	
	signal bitvectord672d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled672d : std_logic := '0';
	signal matchd672d : std_logic := '0';
	
	signal bitvectord673d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled673d : std_logic := '0';
	signal matchd673d : std_logic := '0';
	
	signal bitvectord674d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled674d : std_logic := '0';
	signal matchd674d : std_logic := '0';
	
	signal bitvectord675d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled675d : std_logic := '1';
	signal matchd675d : std_logic := '0';
	
	signal bitvectord676d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled676d : std_logic := '0';
	signal matchd676d : std_logic := '0';
	
	signal bitvectord677d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled677d : std_logic := '0';
	signal matchd677d : std_logic := '0';
	
	signal bitvectord678d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled678d : std_logic := '0';
	signal matchd678d : std_logic := '0';
	
	signal bitvectord679d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled679d : std_logic := '0';
	signal matchd679d : std_logic := '0';
	
	signal bitvectord680d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled680d : std_logic := '0';
	signal matchd680d : std_logic := '0';
	
	signal bitvectord681d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled681d : std_logic := '0';
	signal matchd681d : std_logic := '0';
	
	signal bitvectord682d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled682d : std_logic := '0';
	signal matchd682d : std_logic := '0';
	
	signal bitvectord683d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled683d : std_logic := '0';
	signal matchd683d : std_logic := '0';
	
	signal bitvectord684d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled684d : std_logic := '0';
	signal matchd684d : std_logic := '0';
	
	signal bitvectord685d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled685d : std_logic := '0';
	signal matchd685d : std_logic := '0';
	
	signal bitvectord686d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled686d : std_logic := '0';
	signal matchd686d : std_logic := '0';
	
	signal bitvectord687d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled687d : std_logic := '0';
	signal matchd687d : std_logic := '0';
	
	signal bitvectord688d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled688d : std_logic := '0';
	signal matchd688d : std_logic := '0';
	
	signal bitvectord689d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled689d : std_logic := '0';
	signal matchd689d : std_logic := '0';
	
	signal bitvectord690d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled690d : std_logic := '0';
	signal matchd690d : std_logic := '0';
	
	signal bitvectord691d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled691d : std_logic := '1';
	signal matchd691d : std_logic := '0';
	
	signal bitvectord692d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled692d : std_logic := '0';
	signal matchd692d : std_logic := '0';
	
	signal bitvectord693d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled693d : std_logic := '0';
	signal matchd693d : std_logic := '0';
	
	signal bitvectord694d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled694d : std_logic := '0';
	signal matchd694d : std_logic := '0';
	
	signal bitvectord695d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled695d : std_logic := '0';
	signal matchd695d : std_logic := '0';
	
	signal bitvectord696d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled696d : std_logic := '0';
	signal matchd696d : std_logic := '0';
	
	signal bitvectord697d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled697d : std_logic := '0';
	signal matchd697d : std_logic := '0';
	
	signal bitvectord698d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled698d : std_logic := '0';
	signal matchd698d : std_logic := '0';
	
	signal bitvectord699d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled699d : std_logic := '0';
	signal matchd699d : std_logic := '0';
	
	signal bitvectord700d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled700d : std_logic := '0';
	signal matchd700d : std_logic := '0';
	
	signal bitvectord701d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled701d : std_logic := '0';
	signal matchd701d : std_logic := '0';
	
	signal bitvectord702d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled702d : std_logic := '0';
	signal matchd702d : std_logic := '0';
	
	signal bitvectord703d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled703d : std_logic := '0';
	signal matchd703d : std_logic := '0';
	
	signal bitvectord704d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled704d : std_logic := '0';
	signal matchd704d : std_logic := '0';
	
	signal bitvectord705d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled705d : std_logic := '0';
	signal matchd705d : std_logic := '0';
	
	signal bitvectord706d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled706d : std_logic := '0';
	signal matchd706d : std_logic := '0';
	
	signal bitvectord707d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled707d : std_logic := '0';
	signal matchd707d : std_logic := '0';
	
	signal bitvectord708d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled708d : std_logic := '1';
	signal matchd708d : std_logic := '0';
	
	signal bitvectord709d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled709d : std_logic := '0';
	signal matchd709d : std_logic := '0';
	
	signal bitvectord710d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled710d : std_logic := '0';
	signal matchd710d : std_logic := '0';
	
	signal bitvectord711d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled711d : std_logic := '0';
	signal matchd711d : std_logic := '0';
	
	signal bitvectord712d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled712d : std_logic := '0';
	signal matchd712d : std_logic := '0';
	
	signal bitvectord713d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled713d : std_logic := '0';
	signal matchd713d : std_logic := '0';
	
	signal bitvectord714d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled714d : std_logic := '0';
	signal matchd714d : std_logic := '0';
	
	signal bitvectord715d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled715d : std_logic := '0';
	signal matchd715d : std_logic := '0';
	
	signal bitvectord716d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled716d : std_logic := '0';
	signal matchd716d : std_logic := '0';
	
	signal bitvectord717d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled717d : std_logic := '0';
	signal matchd717d : std_logic := '0';
	
	signal bitvectord718d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled718d : std_logic := '0';
	signal matchd718d : std_logic := '0';
	
	signal bitvectord719d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled719d : std_logic := '0';
	signal matchd719d : std_logic := '0';
	
	signal bitvectord720d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled720d : std_logic := '0';
	signal matchd720d : std_logic := '0';
	
	signal bitvectord721d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled721d : std_logic := '0';
	signal matchd721d : std_logic := '0';
	
	signal bitvectord722d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled722d : std_logic := '0';
	signal matchd722d : std_logic := '0';
	
	signal bitvectord723d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled723d : std_logic := '0';
	signal matchd723d : std_logic := '0';
	
	signal bitvectord724d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled724d : std_logic := '0';
	signal matchd724d : std_logic := '0';
	
	signal bitvectord726d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled726d : std_logic := '1';
	signal matchd726d : std_logic := '0';
	
	signal bitvectord727d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled727d : std_logic := '0';
	signal matchd727d : std_logic := '0';
	
	signal bitvectord728d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled728d : std_logic := '0';
	signal matchd728d : std_logic := '0';
	
	signal bitvectord729d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled729d : std_logic := '0';
	signal matchd729d : std_logic := '0';
	
	signal bitvectord730d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled730d : std_logic := '0';
	signal matchd730d : std_logic := '0';
	
	signal bitvectord731d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled731d : std_logic := '0';
	signal matchd731d : std_logic := '0';
	
	signal bitvectord732d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled732d : std_logic := '0';
	signal matchd732d : std_logic := '0';
	
	signal bitvectord733d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled733d : std_logic := '0';
	signal matchd733d : std_logic := '0';
	
	signal bitvectord734d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled734d : std_logic := '0';
	signal matchd734d : std_logic := '0';
	
	signal bitvectord735d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled735d : std_logic := '0';
	signal matchd735d : std_logic := '0';
	
	signal bitvectord736d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled736d : std_logic := '0';
	signal matchd736d : std_logic := '0';
	
	signal bitvectord737d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled737d : std_logic := '0';
	signal matchd737d : std_logic := '0';
	
	signal bitvectord738d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled738d : std_logic := '0';
	signal matchd738d : std_logic := '0';
	
	signal bitvectord739d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled739d : std_logic := '1';
	signal matchd739d : std_logic := '0';
	
	signal bitvectord740d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled740d : std_logic := '0';
	signal matchd740d : std_logic := '0';
	
	signal bitvectord741d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled741d : std_logic := '0';
	signal matchd741d : std_logic := '0';
	
	signal bitvectord742d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled742d : std_logic := '0';
	signal matchd742d : std_logic := '0';
	
	signal bitvectord743d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled743d : std_logic := '0';
	signal matchd743d : std_logic := '0';
	
	signal bitvectord744d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled744d : std_logic := '0';
	signal matchd744d : std_logic := '0';
	
	signal bitvectord745d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled745d : std_logic := '0';
	signal matchd745d : std_logic := '0';
	
	signal bitvectord746d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled746d : std_logic := '0';
	signal matchd746d : std_logic := '0';
	
	signal bitvectord747d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled747d : std_logic := '0';
	signal matchd747d : std_logic := '0';
	
	signal bitvectord748d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled748d : std_logic := '0';
	signal matchd748d : std_logic := '0';
	
	signal bitvectord749d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled749d : std_logic := '0';
	signal matchd749d : std_logic := '0';
	
	signal bitvectord750d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled750d : std_logic := '0';
	signal matchd750d : std_logic := '0';
	
	signal bitvectord751d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled751d : std_logic := '1';
	signal matchd751d : std_logic := '0';
	
	signal bitvectord752d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled752d : std_logic := '0';
	signal matchd752d : std_logic := '0';
	
	signal bitvectord753d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled753d : std_logic := '0';
	signal matchd753d : std_logic := '0';
	
	signal bitvectord754d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled754d : std_logic := '0';
	signal matchd754d : std_logic := '0';
	
	signal bitvectord755d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled755d : std_logic := '0';
	signal matchd755d : std_logic := '0';
	
	signal bitvectord756d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled756d : std_logic := '0';
	signal matchd756d : std_logic := '0';
	
	signal bitvectord757d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled757d : std_logic := '0';
	signal matchd757d : std_logic := '0';
	
	signal bitvectord758d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled758d : std_logic := '0';
	signal matchd758d : std_logic := '0';
	
	signal bitvectord759d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000";
	signal Enabled759d : std_logic := '0';
	signal matchd759d : std_logic := '0';
	
	signal bitvectord760d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled760d : std_logic := '0';
	signal matchd760d : std_logic := '0';
	
	signal bitvectord761d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled761d : std_logic := '0';
	signal matchd761d : std_logic := '0';
	
	signal bitvectord762d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled762d : std_logic := '0';
	signal matchd762d : std_logic := '0';
	
	signal bitvectord763d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled763d : std_logic := '0';
	signal matchd763d : std_logic := '0';
	
	signal bitvectord764d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled764d : std_logic := '0';
	signal matchd764d : std_logic := '0';
	
	signal bitvectord765d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled765d : std_logic := '0';
	signal matchd765d : std_logic := '0';
	
	signal bitvectord766d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled766d : std_logic := '1';
	signal matchd766d : std_logic := '0';
	
	signal bitvectord767d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled767d : std_logic := '0';
	signal matchd767d : std_logic := '0';
	
	signal bitvectord768d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled768d : std_logic := '0';
	signal matchd768d : std_logic := '0';
	
	signal bitvectord769d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled769d : std_logic := '0';
	signal matchd769d : std_logic := '0';
	
	signal bitvectord770d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled770d : std_logic := '0';
	signal matchd770d : std_logic := '0';
	
	signal bitvectord771d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled771d : std_logic := '0';
	signal matchd771d : std_logic := '0';
	
	signal bitvectord772d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled772d : std_logic := '0';
	signal matchd772d : std_logic := '0';
	
	signal bitvectord773d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled773d : std_logic := '0';
	signal matchd773d : std_logic := '0';
	
	signal bitvectord774d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled774d : std_logic := '0';
	signal matchd774d : std_logic := '0';
	
	signal bitvectord775d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled775d : std_logic := '0';
	signal matchd775d : std_logic := '0';
	
	signal bitvectord776d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled776d : std_logic := '0';
	signal matchd776d : std_logic := '0';
	
	signal bitvectord777d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled777d : std_logic := '1';
	signal matchd777d : std_logic := '0';
	
	signal bitvectord778d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled778d : std_logic := '0';
	signal matchd778d : std_logic := '0';
	
	signal bitvectord779d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled779d : std_logic := '0';
	signal matchd779d : std_logic := '0';
	
	signal bitvectord780d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled780d : std_logic := '0';
	signal matchd780d : std_logic := '0';
	
	signal bitvectord781d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled781d : std_logic := '0';
	signal matchd781d : std_logic := '0';
	
	signal bitvectord782d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled782d : std_logic := '0';
	signal matchd782d : std_logic := '0';
	
	signal bitvectord783d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled783d : std_logic := '0';
	signal matchd783d : std_logic := '0';
	
	signal bitvectord784d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled784d : std_logic := '0';
	signal matchd784d : std_logic := '0';
	
	signal bitvectord785d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled785d : std_logic := '0';
	signal matchd785d : std_logic := '0';
	
	signal bitvectord786d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled786d : std_logic := '0';
	signal matchd786d : std_logic := '0';
	
	signal bitvectord787d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled787d : std_logic := '0';
	signal matchd787d : std_logic := '0';
	
	signal bitvectord788d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled788d : std_logic := '1';
	signal matchd788d : std_logic := '0';
	
	signal bitvectord789d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled789d : std_logic := '0';
	signal matchd789d : std_logic := '0';
	
	signal bitvectord790d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled790d : std_logic := '0';
	signal matchd790d : std_logic := '0';
	
	signal bitvectord791d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled791d : std_logic := '0';
	signal matchd791d : std_logic := '0';
	
	signal bitvectord792d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled792d : std_logic := '0';
	signal matchd792d : std_logic := '0';
	
	signal bitvectord793d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled793d : std_logic := '0';
	signal matchd793d : std_logic := '0';
	
	signal bitvectord794d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled794d : std_logic := '0';
	signal matchd794d : std_logic := '0';
	
	signal bitvectord795d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled795d : std_logic := '0';
	signal matchd795d : std_logic := '0';
	
	signal bitvectord796d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled796d : std_logic := '0';
	signal matchd796d : std_logic := '0';
	
	signal bitvectord797d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled797d : std_logic := '0';
	signal matchd797d : std_logic := '0';
	
	signal bitvectord798d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled798d : std_logic := '0';
	signal matchd798d : std_logic := '0';
	
	signal bitvectord799d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled799d : std_logic := '0';
	signal matchd799d : std_logic := '0';
	
	signal bitvectord800d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled800d : std_logic := '0';
	signal matchd800d : std_logic := '0';
	
	signal bitvectord801d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled801d : std_logic := '0';
	signal matchd801d : std_logic := '0';
	
	signal bitvectord802d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled802d : std_logic := '0';
	signal matchd802d : std_logic := '0';
	
	signal bitvectord803d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled803d : std_logic := '1';
	signal matchd803d : std_logic := '0';
	
	signal bitvectord804d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled804d : std_logic := '0';
	signal matchd804d : std_logic := '0';
	
	signal bitvectord805d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled805d : std_logic := '0';
	signal matchd805d : std_logic := '0';
	
	signal bitvectord806d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled806d : std_logic := '0';
	signal matchd806d : std_logic := '0';
	
	signal bitvectord807d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled807d : std_logic := '0';
	signal matchd807d : std_logic := '0';
	
	signal bitvectord808d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled808d : std_logic := '0';
	signal matchd808d : std_logic := '0';
	
	signal bitvectord809d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled809d : std_logic := '0';
	signal matchd809d : std_logic := '0';
	
	signal bitvectord810d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled810d : std_logic := '0';
	signal matchd810d : std_logic := '0';
	
	signal bitvectord811d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled811d : std_logic := '0';
	signal matchd811d : std_logic := '0';
	
	signal bitvectord812d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled812d : std_logic := '0';
	signal matchd812d : std_logic := '0';
	
	signal bitvectord813d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled813d : std_logic := '0';
	signal matchd813d : std_logic := '0';
	
	signal bitvectord814d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled814d : std_logic := '0';
	signal matchd814d : std_logic := '0';
	
	signal bitvectord815d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled815d : std_logic := '0';
	signal matchd815d : std_logic := '0';
	
	signal bitvectord816d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled816d : std_logic := '0';
	signal matchd816d : std_logic := '0';
	
	signal bitvectord817d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled817d : std_logic := '0';
	signal matchd817d : std_logic := '0';
	
	signal bitvectord819d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled819d : std_logic := '1';
	signal matchd819d : std_logic := '0';
	
	signal bitvectord820d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled820d : std_logic := '0';
	signal matchd820d : std_logic := '0';
	
	signal bitvectord821d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled821d : std_logic := '0';
	signal matchd821d : std_logic := '0';
	
	signal bitvectord822d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled822d : std_logic := '0';
	signal matchd822d : std_logic := '0';
	
	signal bitvectord823d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled823d : std_logic := '0';
	signal matchd823d : std_logic := '0';
	
	signal bitvectord824d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled824d : std_logic := '0';
	signal matchd824d : std_logic := '0';
	
	signal bitvectord825d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled825d : std_logic := '0';
	signal matchd825d : std_logic := '0';
	
	signal bitvectord826d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled826d : std_logic := '0';
	signal matchd826d : std_logic := '0';
	
	signal bitvectord827d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled827d : std_logic := '0';
	signal matchd827d : std_logic := '0';
	
	signal bitvectord828d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled828d : std_logic := '0';
	signal matchd828d : std_logic := '0';
	
	signal bitvectord829d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled829d : std_logic := '0';
	signal matchd829d : std_logic := '0';
	
	signal bitvectord830d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled830d : std_logic := '0';
	signal matchd830d : std_logic := '0';
	
	signal bitvectord831d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled831d : std_logic := '1';
	signal matchd831d : std_logic := '0';
	
	signal bitvectord832d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled832d : std_logic := '0';
	signal matchd832d : std_logic := '0';
	
	signal bitvectord833d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled833d : std_logic := '0';
	signal matchd833d : std_logic := '0';
	
	signal bitvectord834d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled834d : std_logic := '0';
	signal matchd834d : std_logic := '0';
	
	signal bitvectord835d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled835d : std_logic := '0';
	signal matchd835d : std_logic := '0';
	
	signal bitvectord836d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled836d : std_logic := '0';
	signal matchd836d : std_logic := '0';
	
	signal bitvectord837d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled837d : std_logic := '0';
	signal matchd837d : std_logic := '0';
	
	signal bitvectord838d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled838d : std_logic := '0';
	signal matchd838d : std_logic := '0';
	
	signal bitvectord839d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled839d : std_logic := '0';
	signal matchd839d : std_logic := '0';
	
	signal bitvectord840d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000";
	signal Enabled840d : std_logic := '0';
	signal matchd840d : std_logic := '0';
	
	signal bitvectord841d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000";
	signal Enabled841d : std_logic := '0';
	signal matchd841d : std_logic := '0';
	
	signal bitvectord842d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled842d : std_logic := '0';
	signal matchd842d : std_logic := '0';
	
	signal bitvectord843d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled843d : std_logic := '1';
	signal matchd843d : std_logic := '0';
	
	signal bitvectord844d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled844d : std_logic := '0';
	signal matchd844d : std_logic := '0';
	
	signal bitvectord845d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled845d : std_logic := '0';
	signal matchd845d : std_logic := '0';
	
	signal bitvectord846d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled846d : std_logic := '0';
	signal matchd846d : std_logic := '0';
	
	signal bitvectord847d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled847d : std_logic := '0';
	signal matchd847d : std_logic := '0';
	
	signal bitvectord848d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled848d : std_logic := '0';
	signal matchd848d : std_logic := '0';
	
	signal bitvectord849d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled849d : std_logic := '0';
	signal matchd849d : std_logic := '0';
	
	signal bitvectord850d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled850d : std_logic := '0';
	signal matchd850d : std_logic := '0';
	
	signal bitvectord851d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled851d : std_logic := '0';
	signal matchd851d : std_logic := '0';
	
	signal bitvectord852d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled852d : std_logic := '0';
	signal matchd852d : std_logic := '0';
	
	signal bitvectord853d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled853d : std_logic := '0';
	signal matchd853d : std_logic := '0';
	
	signal bitvectord854d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled854d : std_logic := '0';
	signal matchd854d : std_logic := '0';
	
	signal bitvectord855d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled855d : std_logic := '0';
	signal matchd855d : std_logic := '0';
	
	signal bitvectord856d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled856d : std_logic := '0';
	signal matchd856d : std_logic := '0';
	
	signal bitvectord857d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled857d : std_logic := '0';
	signal matchd857d : std_logic := '0';
	
	signal bitvectord858d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled858d : std_logic := '0';
	signal matchd858d : std_logic := '0';
	
	signal bitvectord859d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled859d : std_logic := '0';
	signal matchd859d : std_logic := '0';
	
	signal bitvectord860d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled860d : std_logic := '0';
	signal matchd860d : std_logic := '0';
	
	signal bitvectord861d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled861d : std_logic := '0';
	signal matchd861d : std_logic := '0';
	
	signal bitvectord862d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled862d : std_logic := '0';
	signal matchd862d : std_logic := '0';
	
	signal bitvectord863d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled863d : std_logic := '0';
	signal matchd863d : std_logic := '0';
	
	signal bitvectord864d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled864d : std_logic := '1';
	signal matchd864d : std_logic := '0';
	
	signal bitvectord865d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled865d : std_logic := '0';
	signal matchd865d : std_logic := '0';
	
	signal bitvectord866d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled866d : std_logic := '0';
	signal matchd866d : std_logic := '0';
	
	signal bitvectord867d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled867d : std_logic := '0';
	signal matchd867d : std_logic := '0';
	
	signal bitvectord868d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled868d : std_logic := '0';
	signal matchd868d : std_logic := '0';
	
	signal bitvectord869d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled869d : std_logic := '0';
	signal matchd869d : std_logic := '0';
	
	signal bitvectord870d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled870d : std_logic := '0';
	signal matchd870d : std_logic := '0';
	
	signal bitvectord871d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled871d : std_logic := '0';
	signal matchd871d : std_logic := '0';
	
	signal bitvectord872d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled872d : std_logic := '0';
	signal matchd872d : std_logic := '0';
	
	signal bitvectord873d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled873d : std_logic := '0';
	signal matchd873d : std_logic := '0';
	
	signal bitvectord874d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled874d : std_logic := '0';
	signal matchd874d : std_logic := '0';
	
	signal bitvectord875d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled875d : std_logic := '0';
	signal matchd875d : std_logic := '0';
	
	signal bitvectord876d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled876d : std_logic := '0';
	signal matchd876d : std_logic := '0';
	
	signal bitvectord877d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled877d : std_logic := '0';
	signal matchd877d : std_logic := '0';
	
	signal bitvectord878d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled878d : std_logic := '0';
	signal matchd878d : std_logic := '0';
	
	signal bitvectord879d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled879d : std_logic := '0';
	signal matchd879d : std_logic := '0';
	
	signal bitvectord880d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled880d : std_logic := '0';
	signal matchd880d : std_logic := '0';
	
	signal bitvectord881d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled881d : std_logic := '0';
	signal matchd881d : std_logic := '0';
	
	signal bitvectord882d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled882d : std_logic := '0';
	signal matchd882d : std_logic := '0';
	
	signal bitvectord883d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled883d : std_logic := '0';
	signal matchd883d : std_logic := '0';
	
	signal bitvectord884d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled884d : std_logic := '0';
	signal matchd884d : std_logic := '0';
	
	signal bitvectord885d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled885d : std_logic := '1';
	signal matchd885d : std_logic := '0';
	
	signal bitvectord886d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled886d : std_logic := '0';
	signal matchd886d : std_logic := '0';
	
	signal bitvectord887d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled887d : std_logic := '0';
	signal matchd887d : std_logic := '0';
	
	signal bitvectord888d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled888d : std_logic := '0';
	signal matchd888d : std_logic := '0';
	
	signal bitvectord889d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled889d : std_logic := '0';
	signal matchd889d : std_logic := '0';
	
	signal bitvectord890d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled890d : std_logic := '0';
	signal matchd890d : std_logic := '0';
	
	signal bitvectord891d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled891d : std_logic := '0';
	signal matchd891d : std_logic := '0';
	
	signal bitvectord892d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled892d : std_logic := '0';
	signal matchd892d : std_logic := '0';
	
	signal bitvectord893d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled893d : std_logic := '0';
	signal matchd893d : std_logic := '0';
	
	signal bitvectord894d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled894d : std_logic := '0';
	signal matchd894d : std_logic := '0';
	
	signal bitvectord895d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled895d : std_logic := '0';
	signal matchd895d : std_logic := '0';
	
	signal bitvectord896d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled896d : std_logic := '0';
	signal matchd896d : std_logic := '0';
	
	signal bitvectord897d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled897d : std_logic := '0';
	signal matchd897d : std_logic := '0';
	
	signal bitvectord898d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled898d : std_logic := '0';
	signal matchd898d : std_logic := '0';
	
	signal bitvectord899d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled899d : std_logic := '0';
	signal matchd899d : std_logic := '0';
	
	signal bitvectord900d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled900d : std_logic := '0';
	signal matchd900d : std_logic := '0';
	
	signal bitvectord901d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled901d : std_logic := '0';
	signal matchd901d : std_logic := '0';
	
	signal bitvectord902d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled902d : std_logic := '0';
	signal matchd902d : std_logic := '0';
	
	signal bitvectord903d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled903d : std_logic := '0';
	signal matchd903d : std_logic := '0';
	
	signal bitvectord904d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled904d : std_logic := '0';
	signal matchd904d : std_logic := '0';
	
	signal bitvectord905d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled905d : std_logic := '0';
	signal matchd905d : std_logic := '0';
	
	signal bitvectord907d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled907d : std_logic := '1';
	signal matchd907d : std_logic := '0';
	
	signal bitvectord908d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled908d : std_logic := '0';
	signal matchd908d : std_logic := '0';
	
	signal bitvectord909d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled909d : std_logic := '0';
	signal matchd909d : std_logic := '0';
	
	signal bitvectord910d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled910d : std_logic := '0';
	signal matchd910d : std_logic := '0';
	
	signal bitvectord911d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled911d : std_logic := '0';
	signal matchd911d : std_logic := '0';
	
	signal bitvectord912d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled912d : std_logic := '0';
	signal matchd912d : std_logic := '0';
	
	signal bitvectord913d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled913d : std_logic := '0';
	signal matchd913d : std_logic := '0';
	
	signal bitvectord914d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled914d : std_logic := '0';
	signal matchd914d : std_logic := '0';
	
	signal bitvectord915d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled915d : std_logic := '0';
	signal matchd915d : std_logic := '0';
	
	signal bitvectord916d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled916d : std_logic := '0';
	signal matchd916d : std_logic := '0';
	
	signal bitvectord917d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled917d : std_logic := '0';
	signal matchd917d : std_logic := '0';
	
	signal bitvectord918d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled918d : std_logic := '0';
	signal matchd918d : std_logic := '0';
	
	signal bitvectord919d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled919d : std_logic := '1';
	signal matchd919d : std_logic := '0';
	
	signal bitvectord920d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled920d : std_logic := '0';
	signal matchd920d : std_logic := '0';
	
	signal bitvectord921d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled921d : std_logic := '0';
	signal matchd921d : std_logic := '0';
	
	signal bitvectord922d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled922d : std_logic := '0';
	signal matchd922d : std_logic := '0';
	
	signal bitvectord923d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled923d : std_logic := '0';
	signal matchd923d : std_logic := '0';
	
	signal bitvectord924d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled924d : std_logic := '0';
	signal matchd924d : std_logic := '0';
	
	signal bitvectord925d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled925d : std_logic := '0';
	signal matchd925d : std_logic := '0';
	
	signal bitvectord926d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled926d : std_logic := '0';
	signal matchd926d : std_logic := '0';
	
	signal bitvectord927d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled927d : std_logic := '0';
	signal matchd927d : std_logic := '0';
	
	signal bitvectord928d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled928d : std_logic := '0';
	signal matchd928d : std_logic := '0';
	
	signal bitvectord929d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled929d : std_logic := '0';
	signal matchd929d : std_logic := '0';
	
	signal bitvectord930d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled930d : std_logic := '0';
	signal matchd930d : std_logic := '0';
	
	signal bitvectord931d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled931d : std_logic := '1';
	signal matchd931d : std_logic := '0';
	
	signal bitvectord932d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled932d : std_logic := '0';
	signal matchd932d : std_logic := '0';
	
	signal bitvectord933d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled933d : std_logic := '0';
	signal matchd933d : std_logic := '0';
	
	signal bitvectord934d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled934d : std_logic := '0';
	signal matchd934d : std_logic := '0';
	
	signal bitvectord935d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled935d : std_logic := '0';
	signal matchd935d : std_logic := '0';
	
	signal bitvectord936d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled936d : std_logic := '0';
	signal matchd936d : std_logic := '0';
	
	signal bitvectord937d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled937d : std_logic := '0';
	signal matchd937d : std_logic := '0';
	
	signal bitvectord938d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled938d : std_logic := '0';
	signal matchd938d : std_logic := '0';
	
	signal bitvectord939d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled939d : std_logic := '0';
	signal matchd939d : std_logic := '0';
	
	signal bitvectord940d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled940d : std_logic := '0';
	signal matchd940d : std_logic := '0';
	
	signal bitvectord941d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled941d : std_logic := '0';
	signal matchd941d : std_logic := '0';
	
	signal bitvectord942d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled942d : std_logic := '0';
	signal matchd942d : std_logic := '0';
	
	signal bitvectord943d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled943d : std_logic := '1';
	signal matchd943d : std_logic := '0';
	
	signal bitvectord944d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled944d : std_logic := '0';
	signal matchd944d : std_logic := '0';
	
	signal bitvectord945d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled945d : std_logic := '0';
	signal matchd945d : std_logic := '0';
	
	signal bitvectord946d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled946d : std_logic := '0';
	signal matchd946d : std_logic := '0';
	
	signal bitvectord947d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled947d : std_logic := '0';
	signal matchd947d : std_logic := '0';
	
	signal bitvectord948d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled948d : std_logic := '0';
	signal matchd948d : std_logic := '0';
	
	signal bitvectord949d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled949d : std_logic := '0';
	signal matchd949d : std_logic := '0';
	
	signal bitvectord950d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled950d : std_logic := '0';
	signal matchd950d : std_logic := '0';
	
	signal bitvectord951d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000";
	signal Enabled951d : std_logic := '0';
	signal matchd951d : std_logic := '0';
	
	signal bitvectord952d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled952d : std_logic := '0';
	signal matchd952d : std_logic := '0';
	
	signal bitvectord953d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled953d : std_logic := '0';
	signal matchd953d : std_logic := '0';
	
	signal bitvectord954d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled954d : std_logic := '0';
	signal matchd954d : std_logic := '0';
	
	signal bitvectord955d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111";
	signal Enabled955d : std_logic := '0';
	signal matchd955d : std_logic := '0';
	
	signal bitvectord956d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled956d : std_logic := '0';
	signal matchd956d : std_logic := '0';
	
	signal bitvectord957d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled957d : std_logic := '1';
	signal matchd957d : std_logic := '0';
	
	signal bitvectord958d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled958d : std_logic := '0';
	signal matchd958d : std_logic := '0';
	
	signal bitvectord959d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled959d : std_logic := '0';
	signal matchd959d : std_logic := '0';
	
	signal bitvectord960d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled960d : std_logic := '0';
	signal matchd960d : std_logic := '0';
	
	signal bitvectord961d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled961d : std_logic := '0';
	signal matchd961d : std_logic := '0';
	
	signal bitvectord962d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled962d : std_logic := '0';
	signal matchd962d : std_logic := '0';
	
	signal bitvectord963d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled963d : std_logic := '0';
	signal matchd963d : std_logic := '0';
	
	signal bitvectord964d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled964d : std_logic := '0';
	signal matchd964d : std_logic := '0';
	
	signal bitvectord965d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111";
	signal Enabled965d : std_logic := '0';
	signal matchd965d : std_logic := '0';
	
	signal bitvectord966d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled966d : std_logic := '0';
	signal matchd966d : std_logic := '0';
	
	signal bitvectord967d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled967d : std_logic := '0';
	signal matchd967d : std_logic := '0';
	
	signal bitvectord968d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled968d : std_logic := '0';
	signal matchd968d : std_logic := '0';
	
	signal bitvectord969d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled969d : std_logic := '0';
	signal matchd969d : std_logic := '0';
	
	signal bitvectord970d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled970d : std_logic := '0';
	signal matchd970d : std_logic := '0';
	
	signal bitvectord971d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled971d : std_logic := '1';
	signal matchd971d : std_logic := '0';
	
	signal bitvectord972d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled972d : std_logic := '0';
	signal matchd972d : std_logic := '0';
	
	signal bitvectord973d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled973d : std_logic := '0';
	signal matchd973d : std_logic := '0';
	
	signal bitvectord974d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled974d : std_logic := '0';
	signal matchd974d : std_logic := '0';
	
	signal bitvectord975d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled975d : std_logic := '0';
	signal matchd975d : std_logic := '0';
	
	signal bitvectord976d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled976d : std_logic := '0';
	signal matchd976d : std_logic := '0';
	
	signal bitvectord977d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled977d : std_logic := '0';
	signal matchd977d : std_logic := '0';
	
	signal bitvectord978d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled978d : std_logic := '0';
	signal matchd978d : std_logic := '0';
	
	signal bitvectord979d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled979d : std_logic := '0';
	signal matchd979d : std_logic := '0';
	
	signal bitvectord980d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled980d : std_logic := '0';
	signal matchd980d : std_logic := '0';
	
	signal bitvectord981d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled981d : std_logic := '0';
	signal matchd981d : std_logic := '0';
	
	signal bitvectord982d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled982d : std_logic := '0';
	signal matchd982d : std_logic := '0';
	
	signal bitvectord983d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111";
	signal Enabled983d : std_logic := '0';
	signal matchd983d : std_logic := '0';
	
	signal bitvectord984d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled984d : std_logic := '0';
	signal matchd984d : std_logic := '0';
	
	signal bitvectord986d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled986d : std_logic := '1';
	signal matchd986d : std_logic := '0';
	
	signal bitvectord987d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled987d : std_logic := '0';
	signal matchd987d : std_logic := '0';
	
	signal bitvectord988d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled988d : std_logic := '0';
	signal matchd988d : std_logic := '0';
	
	signal bitvectord989d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled989d : std_logic := '0';
	signal matchd989d : std_logic := '0';
	
	signal bitvectord990d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled990d : std_logic := '0';
	signal matchd990d : std_logic := '0';
	
	signal bitvectord991d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled991d : std_logic := '0';
	signal matchd991d : std_logic := '0';
	
	signal bitvectord992d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled992d : std_logic := '0';
	signal matchd992d : std_logic := '0';
	
	signal bitvectord993d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled993d : std_logic := '0';
	signal matchd993d : std_logic := '0';
	
	signal bitvectord994d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled994d : std_logic := '0';
	signal matchd994d : std_logic := '0';
	
	signal bitvectord995d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled995d : std_logic := '0';
	signal matchd995d : std_logic := '0';
	
	signal bitvectord996d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled996d : std_logic := '0';
	signal matchd996d : std_logic := '0';
	
	signal bitvectord997d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled997d : std_logic := '0';
	signal matchd997d : std_logic := '0';
	
	signal bitvectord998d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled998d : std_logic := '0';
	signal matchd998d : std_logic := '0';
	
	signal bitvectord999d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled999d : std_logic := '0';
	signal matchd999d : std_logic := '0';
	
	signal bitvectord1000d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1000d : std_logic := '0';
	signal matchd1000d : std_logic := '0';
	
	signal bitvectord1001d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1001d : std_logic := '0';
	signal matchd1001d : std_logic := '0';
	
	signal bitvectord1002d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1002d : std_logic := '0';
	signal matchd1002d : std_logic := '0';
	
	signal bitvectord1003d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1003d : std_logic := '0';
	signal matchd1003d : std_logic := '0';
	
	signal bitvectord1004d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1004d : std_logic := '0';
	signal matchd1004d : std_logic := '0';
	
	signal bitvectord1005d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1005d : std_logic := '0';
	signal matchd1005d : std_logic := '0';
	
	signal bitvectord1006d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1006d : std_logic := '0';
	signal matchd1006d : std_logic := '0';
	
	signal bitvectord1007d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1007d : std_logic := '0';
	signal matchd1007d : std_logic := '0';
	
	signal bitvectord1008d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1008d : std_logic := '1';
	signal matchd1008d : std_logic := '0';
	
	signal bitvectord1009d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1009d : std_logic := '0';
	signal matchd1009d : std_logic := '0';
	
	signal bitvectord1010d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1010d : std_logic := '0';
	signal matchd1010d : std_logic := '0';
	
	signal bitvectord1011d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1011d : std_logic := '0';
	signal matchd1011d : std_logic := '0';
	
	signal bitvectord1012d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1012d : std_logic := '0';
	signal matchd1012d : std_logic := '0';
	
	signal bitvectord1013d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1013d : std_logic := '0';
	signal matchd1013d : std_logic := '0';
	
	signal bitvectord1014d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1014d : std_logic := '0';
	signal matchd1014d : std_logic := '0';
	
	signal bitvectord1015d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1015d : std_logic := '0';
	signal matchd1015d : std_logic := '0';
	
	signal bitvectord1016d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1016d : std_logic := '0';
	signal matchd1016d : std_logic := '0';
	
	signal bitvectord1017d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1017d : std_logic := '0';
	signal matchd1017d : std_logic := '0';
	
	signal bitvectord1018d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1018d : std_logic := '0';
	signal matchd1018d : std_logic := '0';
	
	signal bitvectord1019d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1019d : std_logic := '0';
	signal matchd1019d : std_logic := '0';
	
	signal bitvectord1020d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1020d : std_logic := '0';
	signal matchd1020d : std_logic := '0';
	
	signal bitvectord1021d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1021d : std_logic := '0';
	signal matchd1021d : std_logic := '0';
	
	signal bitvectord1022d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1022d : std_logic := '0';
	signal matchd1022d : std_logic := '0';
	
	signal bitvectord1023d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1023d : std_logic := '0';
	signal matchd1023d : std_logic := '0';
	
	signal bitvectord1024d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1024d : std_logic := '0';
	signal matchd1024d : std_logic := '0';
	
	signal bitvectord1025d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1025d : std_logic := '0';
	signal matchd1025d : std_logic := '0';
	
	signal bitvectord1026d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1026d : std_logic := '0';
	signal matchd1026d : std_logic := '0';
	
	signal bitvectord1027d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1027d : std_logic := '0';
	signal matchd1027d : std_logic := '0';
	
	signal bitvectord1028d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1028d : std_logic := '0';
	signal matchd1028d : std_logic := '0';
	
	signal bitvectord1029d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1029d : std_logic := '1';
	signal matchd1029d : std_logic := '0';
	
	signal bitvectord1030d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1030d : std_logic := '0';
	signal matchd1030d : std_logic := '0';
	
	signal bitvectord1031d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1031d : std_logic := '0';
	signal matchd1031d : std_logic := '0';
	
	signal bitvectord1032d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1032d : std_logic := '0';
	signal matchd1032d : std_logic := '0';
	
	signal bitvectord1033d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1033d : std_logic := '0';
	signal matchd1033d : std_logic := '0';
	
	signal bitvectord1034d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1034d : std_logic := '0';
	signal matchd1034d : std_logic := '0';
	
	signal bitvectord1035d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1035d : std_logic := '0';
	signal matchd1035d : std_logic := '0';
	
	signal bitvectord1036d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1036d : std_logic := '0';
	signal matchd1036d : std_logic := '0';
	
	signal bitvectord1037d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1037d : std_logic := '0';
	signal matchd1037d : std_logic := '0';
	
	signal bitvectord1038d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1038d : std_logic := '0';
	signal matchd1038d : std_logic := '0';
	
	signal bitvectord1039d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1039d : std_logic := '0';
	signal matchd1039d : std_logic := '0';
	
	signal bitvectord1040d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1040d : std_logic := '1';
	signal matchd1040d : std_logic := '0';
	
	signal bitvectord1041d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1041d : std_logic := '0';
	signal matchd1041d : std_logic := '0';
	
	signal bitvectord1042d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1042d : std_logic := '0';
	signal matchd1042d : std_logic := '0';
	
	signal bitvectord1043d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1043d : std_logic := '0';
	signal matchd1043d : std_logic := '0';
	
	signal bitvectord1044d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1044d : std_logic := '0';
	signal matchd1044d : std_logic := '0';
	
	signal bitvectord1045d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1045d : std_logic := '0';
	signal matchd1045d : std_logic := '0';
	
	signal bitvectord1046d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1046d : std_logic := '0';
	signal matchd1046d : std_logic := '0';
	
	signal bitvectord1047d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1047d : std_logic := '0';
	signal matchd1047d : std_logic := '0';
	
	signal bitvectord1048d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1048d : std_logic := '0';
	signal matchd1048d : std_logic := '0';
	
	signal bitvectord1049d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1049d : std_logic := '0';
	signal matchd1049d : std_logic := '0';
	
	signal bitvectord1050d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1050d : std_logic := '0';
	signal matchd1050d : std_logic := '0';
	
	signal bitvectord1051d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1051d : std_logic := '0';
	signal matchd1051d : std_logic := '0';
	
	signal bitvectord1052d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1052d : std_logic := '1';
	signal matchd1052d : std_logic := '0';
	
	signal bitvectord1053d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1053d : std_logic := '0';
	signal matchd1053d : std_logic := '0';
	
	signal bitvectord1054d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1054d : std_logic := '0';
	signal matchd1054d : std_logic := '0';
	
	signal bitvectord1055d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1055d : std_logic := '0';
	signal matchd1055d : std_logic := '0';
	
	signal bitvectord1056d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1056d : std_logic := '0';
	signal matchd1056d : std_logic := '0';
	
	signal bitvectord1057d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1057d : std_logic := '0';
	signal matchd1057d : std_logic := '0';
	
	signal bitvectord1058d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1058d : std_logic := '0';
	signal matchd1058d : std_logic := '0';
	
	signal bitvectord1059d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1059d : std_logic := '0';
	signal matchd1059d : std_logic := '0';
	
	signal bitvectord1060d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1060d : std_logic := '0';
	signal matchd1060d : std_logic := '0';
	
	signal bitvectord1061d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1061d : std_logic := '0';
	signal matchd1061d : std_logic := '0';
	
	signal bitvectord1062d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1062d : std_logic := '0';
	signal matchd1062d : std_logic := '0';
	
	signal bitvectord1063d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1063d : std_logic := '0';
	signal matchd1063d : std_logic := '0';
	
	signal bitvectord1064d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1064d : std_logic := '1';
	signal matchd1064d : std_logic := '0';
	
	signal bitvectord1065d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1065d : std_logic := '0';
	signal matchd1065d : std_logic := '0';
	
	signal bitvectord1066d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1066d : std_logic := '0';
	signal matchd1066d : std_logic := '0';
	
	signal bitvectord1067d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1067d : std_logic := '0';
	signal matchd1067d : std_logic := '0';
	
	signal bitvectord1068d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1068d : std_logic := '0';
	signal matchd1068d : std_logic := '0';
	
	signal bitvectord1069d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1069d : std_logic := '0';
	signal matchd1069d : std_logic := '0';
	
	signal bitvectord1070d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1070d : std_logic := '0';
	signal matchd1070d : std_logic := '0';
	
	signal bitvectord1071d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1071d : std_logic := '0';
	signal matchd1071d : std_logic := '0';
	
	signal bitvectord1072d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1072d : std_logic := '0';
	signal matchd1072d : std_logic := '0';
	
	signal bitvectord1073d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1073d : std_logic := '0';
	signal matchd1073d : std_logic := '0';
	
	signal bitvectord1074d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1074d : std_logic := '0';
	signal matchd1074d : std_logic := '0';
	
	signal bitvectord1075d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1075d : std_logic := '0';
	signal matchd1075d : std_logic := '0';
	
	signal bitvectord1076d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1076d : std_logic := '1';
	signal matchd1076d : std_logic := '0';
	
	signal bitvectord1077d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1077d : std_logic := '0';
	signal matchd1077d : std_logic := '0';
	
	signal bitvectord1078d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1078d : std_logic := '0';
	signal matchd1078d : std_logic := '0';
	
	signal bitvectord1079d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1079d : std_logic := '0';
	signal matchd1079d : std_logic := '0';
	
	signal bitvectord1080d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1080d : std_logic := '0';
	signal matchd1080d : std_logic := '0';
	
	signal bitvectord1081d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1081d : std_logic := '0';
	signal matchd1081d : std_logic := '0';
	
	signal bitvectord1082d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1082d : std_logic := '0';
	signal matchd1082d : std_logic := '0';
	
	signal bitvectord1083d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1083d : std_logic := '0';
	signal matchd1083d : std_logic := '0';
	
	signal bitvectord1084d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1084d : std_logic := '0';
	signal matchd1084d : std_logic := '0';
	
	signal bitvectord1085d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1085d : std_logic := '1';
	signal matchd1085d : std_logic := '0';
	
	signal bitvectord1086d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1086d : std_logic := '0';
	signal matchd1086d : std_logic := '0';
	
	signal bitvectord1087d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1087d : std_logic := '0';
	signal matchd1087d : std_logic := '0';
	
	signal bitvectord1088d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled1088d : std_logic := '0';
	signal matchd1088d : std_logic := '0';
	
	signal bitvectord1089d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1089d : std_logic := '0';
	signal matchd1089d : std_logic := '0';
	
	signal bitvectord1090d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1090d : std_logic := '0';
	signal matchd1090d : std_logic := '0';
	
	signal bitvectord1091d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1091d : std_logic := '0';
	signal matchd1091d : std_logic := '0';
	
	signal bitvectord1092d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1092d : std_logic := '0';
	signal matchd1092d : std_logic := '0';
	
	signal bitvectord1093d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1093d : std_logic := '0';
	signal matchd1093d : std_logic := '0';
	
	signal bitvectord1094d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1094d : std_logic := '0';
	signal matchd1094d : std_logic := '0';
	
	signal bitvectord1095d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1095d : std_logic := '0';
	signal matchd1095d : std_logic := '0';
	
	signal bitvectord1096d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1096d : std_logic := '0';
	signal matchd1096d : std_logic := '0';
	
	signal bitvectord1097d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1097d : std_logic := '0';
	signal matchd1097d : std_logic := '0';
	
	signal bitvectord1098d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1098d : std_logic := '0';
	signal matchd1098d : std_logic := '0';
	
	signal bitvectord1099d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1099d : std_logic := '0';
	signal matchd1099d : std_logic := '0';
	
	signal bitvectord1100d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1100d : std_logic := '0';
	signal matchd1100d : std_logic := '0';
	
	signal bitvectord1101d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1101d : std_logic := '0';
	signal matchd1101d : std_logic := '0';
	
	signal bitvectord1102d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1102d : std_logic := '1';
	signal matchd1102d : std_logic := '0';
	
	signal bitvectord1103d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1103d : std_logic := '0';
	signal matchd1103d : std_logic := '0';
	
	signal bitvectord1104d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1104d : std_logic := '0';
	signal matchd1104d : std_logic := '0';
	
	signal bitvectord1105d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1105d : std_logic := '0';
	signal matchd1105d : std_logic := '0';
	
	signal bitvectord1106d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1106d : std_logic := '0';
	signal matchd1106d : std_logic := '0';
	
	signal bitvectord1107d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1107d : std_logic := '0';
	signal matchd1107d : std_logic := '0';
	
	signal bitvectord1108d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1108d : std_logic := '0';
	signal matchd1108d : std_logic := '0';
	
	signal bitvectord1109d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1109d : std_logic := '0';
	signal matchd1109d : std_logic := '0';
	
	signal bitvectord1110d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1110d : std_logic := '0';
	signal matchd1110d : std_logic := '0';
	
	signal bitvectord1111d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled1111d : std_logic := '0';
	signal matchd1111d : std_logic := '0';
	
	signal bitvectord1112d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1112d : std_logic := '0';
	signal matchd1112d : std_logic := '0';
	
	signal bitvectord1113d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1113d : std_logic := '0';
	signal matchd1113d : std_logic := '0';
	
	signal bitvectord1114d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1114d : std_logic := '0';
	signal matchd1114d : std_logic := '0';
	
	signal bitvectord1115d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1115d : std_logic := '0';
	signal matchd1115d : std_logic := '0';
	
	signal bitvectord1116d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1116d : std_logic := '0';
	signal matchd1116d : std_logic := '0';
	
	signal bitvectord1117d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1117d : std_logic := '0';
	signal matchd1117d : std_logic := '0';
	
	signal bitvectord1118d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1118d : std_logic := '0';
	signal matchd1118d : std_logic := '0';
	
	signal bitvectord1120d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1120d : std_logic := '1';
	signal matchd1120d : std_logic := '0';
	
	signal bitvectord1121d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1121d : std_logic := '0';
	signal matchd1121d : std_logic := '0';
	
	signal bitvectord1122d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1122d : std_logic := '0';
	signal matchd1122d : std_logic := '0';
	
	signal bitvectord1123d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1123d : std_logic := '0';
	signal matchd1123d : std_logic := '0';
	
	signal bitvectord1124d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1124d : std_logic := '0';
	signal matchd1124d : std_logic := '0';
	
	signal bitvectord1125d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1125d : std_logic := '0';
	signal matchd1125d : std_logic := '0';
	
	signal bitvectord1126d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1126d : std_logic := '0';
	signal matchd1126d : std_logic := '0';
	
	signal bitvectord1127d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1127d : std_logic := '0';
	signal matchd1127d : std_logic := '0';
	
	signal bitvectord1128d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1128d : std_logic := '0';
	signal matchd1128d : std_logic := '0';
	
	signal bitvectord1129d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1129d : std_logic := '0';
	signal matchd1129d : std_logic := '0';
	
	signal bitvectord1130d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1130d : std_logic := '0';
	signal matchd1130d : std_logic := '0';
	
	signal bitvectord1131d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1131d : std_logic := '1';
	signal matchd1131d : std_logic := '0';
	
	signal bitvectord1132d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1132d : std_logic := '0';
	signal matchd1132d : std_logic := '0';
	
	signal bitvectord1133d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1133d : std_logic := '0';
	signal matchd1133d : std_logic := '0';
	
	signal bitvectord1134d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1134d : std_logic := '0';
	signal matchd1134d : std_logic := '0';
	
	signal bitvectord1135d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1135d : std_logic := '0';
	signal matchd1135d : std_logic := '0';
	
	signal bitvectord1136d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1136d : std_logic := '0';
	signal matchd1136d : std_logic := '0';
	
	signal bitvectord1137d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1137d : std_logic := '0';
	signal matchd1137d : std_logic := '0';
	
	signal bitvectord1138d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1138d : std_logic := '0';
	signal matchd1138d : std_logic := '0';
	
	signal bitvectord1139d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1139d : std_logic := '0';
	signal matchd1139d : std_logic := '0';
	
	signal bitvectord1140d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1140d : std_logic := '0';
	signal matchd1140d : std_logic := '0';
	
	signal bitvectord1141d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1141d : std_logic := '0';
	signal matchd1141d : std_logic := '0';
	
	signal bitvectord1142d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1142d : std_logic := '0';
	signal matchd1142d : std_logic := '0';
	
	signal bitvectord1143d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1143d : std_logic := '1';
	signal matchd1143d : std_logic := '0';
	
	signal bitvectord1144d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1144d : std_logic := '0';
	signal matchd1144d : std_logic := '0';
	
	signal bitvectord1145d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1145d : std_logic := '0';
	signal matchd1145d : std_logic := '0';
	
	signal bitvectord1146d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1146d : std_logic := '0';
	signal matchd1146d : std_logic := '0';
	
	signal bitvectord1147d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1147d : std_logic := '0';
	signal matchd1147d : std_logic := '0';
	
	signal bitvectord1148d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1148d : std_logic := '0';
	signal matchd1148d : std_logic := '0';
	
	signal bitvectord1149d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1149d : std_logic := '0';
	signal matchd1149d : std_logic := '0';
	
	signal bitvectord1150d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1150d : std_logic := '0';
	signal matchd1150d : std_logic := '0';
	
	signal bitvectord1151d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1151d : std_logic := '0';
	signal matchd1151d : std_logic := '0';
	
	signal bitvectord1152d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1152d : std_logic := '0';
	signal matchd1152d : std_logic := '0';
	
	signal bitvectord1153d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1153d : std_logic := '1';
	signal matchd1153d : std_logic := '0';
	
	signal bitvectord1154d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1154d : std_logic := '0';
	signal matchd1154d : std_logic := '0';
	
	signal bitvectord1155d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1155d : std_logic := '0';
	signal matchd1155d : std_logic := '0';
	
	signal bitvectord1156d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1156d : std_logic := '0';
	signal matchd1156d : std_logic := '0';
	
	signal bitvectord1157d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1157d : std_logic := '0';
	signal matchd1157d : std_logic := '0';
	
	signal bitvectord1158d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1158d : std_logic := '0';
	signal matchd1158d : std_logic := '0';
	
	signal bitvectord1159d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1159d : std_logic := '0';
	signal matchd1159d : std_logic := '0';
	
	signal bitvectord1160d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1160d : std_logic := '0';
	signal matchd1160d : std_logic := '0';
	
	signal bitvectord1161d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled1161d : std_logic := '0';
	signal matchd1161d : std_logic := '0';
	
	signal bitvectord1162d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1162d : std_logic := '0';
	signal matchd1162d : std_logic := '0';
	
	signal bitvectord1163d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1163d : std_logic := '0';
	signal matchd1163d : std_logic := '0';
	
	signal bitvectord1164d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1164d : std_logic := '0';
	signal matchd1164d : std_logic := '0';
	
	signal bitvectord1165d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1165d : std_logic := '0';
	signal matchd1165d : std_logic := '0';
	
	signal bitvectord1166d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1166d : std_logic := '0';
	signal matchd1166d : std_logic := '0';
	
	signal bitvectord1167d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1167d : std_logic := '0';
	signal matchd1167d : std_logic := '0';
	
	signal bitvectord1168d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1168d : std_logic := '0';
	signal matchd1168d : std_logic := '0';
	
	signal bitvectord1169d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1169d : std_logic := '1';
	signal matchd1169d : std_logic := '0';
	
	signal bitvectord1170d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1170d : std_logic := '0';
	signal matchd1170d : std_logic := '0';
	
	signal bitvectord1171d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1171d : std_logic := '0';
	signal matchd1171d : std_logic := '0';
	
	signal bitvectord1172d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1172d : std_logic := '0';
	signal matchd1172d : std_logic := '0';
	
	signal bitvectord1173d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1173d : std_logic := '0';
	signal matchd1173d : std_logic := '0';
	
	signal bitvectord1174d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1174d : std_logic := '0';
	signal matchd1174d : std_logic := '0';
	
	signal bitvectord1175d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1175d : std_logic := '0';
	signal matchd1175d : std_logic := '0';
	
	signal bitvectord1176d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1176d : std_logic := '0';
	signal matchd1176d : std_logic := '0';
	
	signal bitvectord1177d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1177d : std_logic := '0';
	signal matchd1177d : std_logic := '0';
	
	signal bitvectord1178d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1178d : std_logic := '0';
	signal matchd1178d : std_logic := '0';
	
	signal bitvectord1179d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1179d : std_logic := '0';
	signal matchd1179d : std_logic := '0';
	
	signal bitvectord1180d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1180d : std_logic := '0';
	signal matchd1180d : std_logic := '0';
	
	signal bitvectord1181d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1181d : std_logic := '0';
	signal matchd1181d : std_logic := '0';
	
	signal bitvectord1182d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1182d : std_logic := '1';
	signal matchd1182d : std_logic := '0';
	
	signal bitvectord1183d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1183d : std_logic := '0';
	signal matchd1183d : std_logic := '0';
	
	signal bitvectord1184d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1184d : std_logic := '0';
	signal matchd1184d : std_logic := '0';
	
	signal bitvectord1185d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1185d : std_logic := '0';
	signal matchd1185d : std_logic := '0';
	
	signal bitvectord1186d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1186d : std_logic := '0';
	signal matchd1186d : std_logic := '0';
	
	signal bitvectord1187d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1187d : std_logic := '0';
	signal matchd1187d : std_logic := '0';
	
	signal bitvectord1188d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1188d : std_logic := '0';
	signal matchd1188d : std_logic := '0';
	
	signal bitvectord1189d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1189d : std_logic := '0';
	signal matchd1189d : std_logic := '0';
	
	signal bitvectord1190d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1190d : std_logic := '0';
	signal matchd1190d : std_logic := '0';
	
	signal bitvectord1191d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1191d : std_logic := '0';
	signal matchd1191d : std_logic := '0';
	
	signal bitvectord1192d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1192d : std_logic := '0';
	signal matchd1192d : std_logic := '0';
	
	signal bitvectord1193d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1193d : std_logic := '1';
	signal matchd1193d : std_logic := '0';
	
	signal bitvectord1194d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1194d : std_logic := '0';
	signal matchd1194d : std_logic := '0';
	
	signal bitvectord1195d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1195d : std_logic := '0';
	signal matchd1195d : std_logic := '0';
	
	signal bitvectord1196d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1196d : std_logic := '0';
	signal matchd1196d : std_logic := '0';
	
	signal bitvectord1197d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1197d : std_logic := '0';
	signal matchd1197d : std_logic := '0';
	
	signal bitvectord1198d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1198d : std_logic := '0';
	signal matchd1198d : std_logic := '0';
	
	signal bitvectord1199d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1199d : std_logic := '0';
	signal matchd1199d : std_logic := '0';
	
	signal bitvectord1200d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1200d : std_logic := '0';
	signal matchd1200d : std_logic := '0';
	
	signal bitvectord1201d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1201d : std_logic := '0';
	signal matchd1201d : std_logic := '0';
	
	signal bitvectord1202d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1202d : std_logic := '0';
	signal matchd1202d : std_logic := '0';
	
	signal bitvectord1203d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1203d : std_logic := '0';
	signal matchd1203d : std_logic := '0';
	
	signal bitvectord1204d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1204d : std_logic := '0';
	signal matchd1204d : std_logic := '0';
	
	signal bitvectord1205d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1205d : std_logic := '0';
	signal matchd1205d : std_logic := '0';
	
	signal bitvectord1206d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1206d : std_logic := '0';
	signal matchd1206d : std_logic := '0';
	
	signal bitvectord1207d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1207d : std_logic := '0';
	signal matchd1207d : std_logic := '0';
	
	signal bitvectord1208d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1208d : std_logic := '0';
	signal matchd1208d : std_logic := '0';
	
	signal bitvectord1209d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1209d : std_logic := '0';
	signal matchd1209d : std_logic := '0';
	
	signal bitvectord1210d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1210d : std_logic := '0';
	signal matchd1210d : std_logic := '0';
	
	signal bitvectord1211d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1211d : std_logic := '0';
	signal matchd1211d : std_logic := '0';
	
	signal bitvectord1212d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1212d : std_logic := '0';
	signal matchd1212d : std_logic := '0';
	
	signal bitvectord1213d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1213d : std_logic := '0';
	signal matchd1213d : std_logic := '0';
	
	signal bitvectord1214d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1214d : std_logic := '1';
	signal matchd1214d : std_logic := '0';
	
	signal bitvectord1215d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1215d : std_logic := '0';
	signal matchd1215d : std_logic := '0';
	
	signal bitvectord1216d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1216d : std_logic := '0';
	signal matchd1216d : std_logic := '0';
	
	signal bitvectord1217d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1217d : std_logic := '0';
	signal matchd1217d : std_logic := '0';
	
	signal bitvectord1218d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1218d : std_logic := '0';
	signal matchd1218d : std_logic := '0';
	
	signal bitvectord1219d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1219d : std_logic := '0';
	signal matchd1219d : std_logic := '0';
	
	signal bitvectord1220d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1220d : std_logic := '0';
	signal matchd1220d : std_logic := '0';
	
	signal bitvectord1221d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1221d : std_logic := '0';
	signal matchd1221d : std_logic := '0';
	
	signal bitvectord1222d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1222d : std_logic := '0';
	signal matchd1222d : std_logic := '0';
	
	signal bitvectord1223d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1223d : std_logic := '0';
	signal matchd1223d : std_logic := '0';
	
	signal bitvectord1224d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1224d : std_logic := '0';
	signal matchd1224d : std_logic := '0';
	
	signal bitvectord1225d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1225d : std_logic := '1';
	signal matchd1225d : std_logic := '0';
	
	signal bitvectord1226d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1226d : std_logic := '0';
	signal matchd1226d : std_logic := '0';
	
	signal bitvectord1227d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1227d : std_logic := '0';
	signal matchd1227d : std_logic := '0';
	
	signal bitvectord1228d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1228d : std_logic := '0';
	signal matchd1228d : std_logic := '0';
	
	signal bitvectord1229d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1229d : std_logic := '0';
	signal matchd1229d : std_logic := '0';
	
	signal bitvectord1230d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1230d : std_logic := '0';
	signal matchd1230d : std_logic := '0';
	
	signal bitvectord1231d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1231d : std_logic := '0';
	signal matchd1231d : std_logic := '0';
	
	signal bitvectord1232d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1232d : std_logic := '0';
	signal matchd1232d : std_logic := '0';
	
	signal bitvectord1233d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1233d : std_logic := '0';
	signal matchd1233d : std_logic := '0';
	
	signal bitvectord1234d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1234d : std_logic := '0';
	signal matchd1234d : std_logic := '0';
	
	signal bitvectord1235d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1235d : std_logic := '0';
	signal matchd1235d : std_logic := '0';
	
	signal bitvectord1236d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1236d : std_logic := '0';
	signal matchd1236d : std_logic := '0';
	
	signal bitvectord1237d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1237d : std_logic := '0';
	signal matchd1237d : std_logic := '0';
	
	signal bitvectord1238d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1238d : std_logic := '0';
	signal matchd1238d : std_logic := '0';
	
	signal bitvectord1239d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1239d : std_logic := '0';
	signal matchd1239d : std_logic := '0';
	
	signal bitvectord1240d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1240d : std_logic := '0';
	signal matchd1240d : std_logic := '0';
	
	signal bitvectord1241d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1241d : std_logic := '0';
	signal matchd1241d : std_logic := '0';
	
	signal bitvectord1242d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1242d : std_logic := '1';
	signal matchd1242d : std_logic := '0';
	
	signal bitvectord1243d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1243d : std_logic := '0';
	signal matchd1243d : std_logic := '0';
	
	signal bitvectord1244d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1244d : std_logic := '0';
	signal matchd1244d : std_logic := '0';
	
	signal bitvectord1245d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1245d : std_logic := '0';
	signal matchd1245d : std_logic := '0';
	
	signal bitvectord1246d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1246d : std_logic := '0';
	signal matchd1246d : std_logic := '0';
	
	signal bitvectord1247d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1247d : std_logic := '0';
	signal matchd1247d : std_logic := '0';
	
	signal bitvectord1248d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1248d : std_logic := '0';
	signal matchd1248d : std_logic := '0';
	
	signal bitvectord1249d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1249d : std_logic := '0';
	signal matchd1249d : std_logic := '0';
	
	signal bitvectord1250d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1250d : std_logic := '0';
	signal matchd1250d : std_logic := '0';
	
	signal bitvectord1251d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1251d : std_logic := '0';
	signal matchd1251d : std_logic := '0';
	
	signal bitvectord1252d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1252d : std_logic := '0';
	signal matchd1252d : std_logic := '0';
	
	signal bitvectord1253d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1253d : std_logic := '0';
	signal matchd1253d : std_logic := '0';
	
	signal bitvectord1254d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1254d : std_logic := '1';
	signal matchd1254d : std_logic := '0';
	
	signal bitvectord1255d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1255d : std_logic := '0';
	signal matchd1255d : std_logic := '0';
	
	signal bitvectord1256d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1256d : std_logic := '0';
	signal matchd1256d : std_logic := '0';
	
	signal bitvectord1257d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1257d : std_logic := '0';
	signal matchd1257d : std_logic := '0';
	
	signal bitvectord1258d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1258d : std_logic := '0';
	signal matchd1258d : std_logic := '0';
	
	signal bitvectord1259d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1259d : std_logic := '0';
	signal matchd1259d : std_logic := '0';
	
	signal bitvectord1260d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1260d : std_logic := '0';
	signal matchd1260d : std_logic := '0';
	
	signal bitvectord1261d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1261d : std_logic := '0';
	signal matchd1261d : std_logic := '0';
	
	signal bitvectord1262d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1262d : std_logic := '0';
	signal matchd1262d : std_logic := '0';
	
	signal bitvectord1263d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1263d : std_logic := '0';
	signal matchd1263d : std_logic := '0';
	
	signal bitvectord1264d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1264d : std_logic := '0';
	signal matchd1264d : std_logic := '0';
	
	signal bitvectord1265d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1265d : std_logic := '0';
	signal matchd1265d : std_logic := '0';
	
	signal bitvectord1266d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1266d : std_logic := '0';
	signal matchd1266d : std_logic := '0';
	
	signal bitvectord1267d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1267d : std_logic := '1';
	signal matchd1267d : std_logic := '0';
	
	signal bitvectord1268d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1268d : std_logic := '0';
	signal matchd1268d : std_logic := '0';
	
	signal bitvectord1269d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1269d : std_logic := '0';
	signal matchd1269d : std_logic := '0';
	
	signal bitvectord1270d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled1270d : std_logic := '0';
	signal matchd1270d : std_logic := '0';
	
	signal bitvectord1271d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1271d : std_logic := '0';
	signal matchd1271d : std_logic := '0';
	
	signal bitvectord1272d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1272d : std_logic := '0';
	signal matchd1272d : std_logic := '0';
	
	signal bitvectord1273d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1273d : std_logic := '0';
	signal matchd1273d : std_logic := '0';
	
	signal bitvectord1274d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1274d : std_logic := '0';
	signal matchd1274d : std_logic := '0';
	
	signal bitvectord1275d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1275d : std_logic := '0';
	signal matchd1275d : std_logic := '0';
	
	signal bitvectord1276d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1276d : std_logic := '0';
	signal matchd1276d : std_logic := '0';
	
	signal bitvectord1277d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1277d : std_logic := '0';
	signal matchd1277d : std_logic := '0';
	
	signal bitvectord1278d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1278d : std_logic := '0';
	signal matchd1278d : std_logic := '0';
	
	signal bitvectord1279d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1279d : std_logic := '0';
	signal matchd1279d : std_logic := '0';
	
	signal bitvectord1280d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000";
	signal Enabled1280d : std_logic := '0';
	signal matchd1280d : std_logic := '0';
	
	signal bitvectord1281d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000";
	signal Enabled1281d : std_logic := '0';
	signal matchd1281d : std_logic := '0';
	
	signal bitvectord1282d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1282d : std_logic := '0';
	signal matchd1282d : std_logic := '0';
	
	signal bitvectord1283d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1283d : std_logic := '1';
	signal matchd1283d : std_logic := '0';
	
	signal bitvectord1284d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1284d : std_logic := '0';
	signal matchd1284d : std_logic := '0';
	
	signal bitvectord1285d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1285d : std_logic := '0';
	signal matchd1285d : std_logic := '0';
	
	signal bitvectord1286d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1286d : std_logic := '0';
	signal matchd1286d : std_logic := '0';
	
	signal bitvectord1287d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1287d : std_logic := '0';
	signal matchd1287d : std_logic := '0';
	
	signal bitvectord1288d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1288d : std_logic := '0';
	signal matchd1288d : std_logic := '0';
	
	signal bitvectord1289d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1289d : std_logic := '0';
	signal matchd1289d : std_logic := '0';
	
	signal bitvectord1290d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1290d : std_logic := '0';
	signal matchd1290d : std_logic := '0';
	
	signal bitvectord1291d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1291d : std_logic := '0';
	signal matchd1291d : std_logic := '0';
	
	signal bitvectord1292d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled1292d : std_logic := '0';
	signal matchd1292d : std_logic := '0';
	
	signal bitvectord1293d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1293d : std_logic := '0';
	signal matchd1293d : std_logic := '0';
	
	signal bitvectord1294d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1294d : std_logic := '0';
	signal matchd1294d : std_logic := '0';
	
	signal bitvectord1295d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1295d : std_logic := '0';
	signal matchd1295d : std_logic := '0';
	
	signal bitvectord1296d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000";
	signal Enabled1296d : std_logic := '0';
	signal matchd1296d : std_logic := '0';
	
	signal bitvectord1297d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000";
	signal Enabled1297d : std_logic := '0';
	signal matchd1297d : std_logic := '0';
	
	signal bitvectord1298d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1298d : std_logic := '0';
	signal matchd1298d : std_logic := '0';
	
	signal bitvectord1300d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1300d : std_logic := '1';
	signal matchd1300d : std_logic := '0';
	
	signal bitvectord1301d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1301d : std_logic := '0';
	signal matchd1301d : std_logic := '0';
	
	signal bitvectord1302d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1302d : std_logic := '0';
	signal matchd1302d : std_logic := '0';
	
	signal bitvectord1303d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1303d : std_logic := '0';
	signal matchd1303d : std_logic := '0';
	
	signal bitvectord1304d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1304d : std_logic := '0';
	signal matchd1304d : std_logic := '0';
	
	signal bitvectord1305d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled1305d : std_logic := '0';
	signal matchd1305d : std_logic := '0';
	
	signal bitvectord1306d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1306d : std_logic := '0';
	signal matchd1306d : std_logic := '0';
	
	signal bitvectord1307d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1307d : std_logic := '0';
	signal matchd1307d : std_logic := '0';
	
	signal bitvectord1308d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1308d : std_logic := '0';
	signal matchd1308d : std_logic := '0';
	
	signal bitvectord1309d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1309d : std_logic := '0';
	signal matchd1309d : std_logic := '0';
	
	signal bitvectord1310d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1310d : std_logic := '0';
	signal matchd1310d : std_logic := '0';
	
	signal bitvectord1311d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1311d : std_logic := '0';
	signal matchd1311d : std_logic := '0';
	
	signal bitvectord1312d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1312d : std_logic := '0';
	signal matchd1312d : std_logic := '0';
	
	signal bitvectord1313d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1313d : std_logic := '1';
	signal matchd1313d : std_logic := '0';
	
	signal bitvectord1314d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1314d : std_logic := '0';
	signal matchd1314d : std_logic := '0';
	
	signal bitvectord1315d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1315d : std_logic := '0';
	signal matchd1315d : std_logic := '0';
	
	signal bitvectord1316d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1316d : std_logic := '0';
	signal matchd1316d : std_logic := '0';
	
	signal bitvectord1317d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1317d : std_logic := '0';
	signal matchd1317d : std_logic := '0';
	
	signal bitvectord1318d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1318d : std_logic := '0';
	signal matchd1318d : std_logic := '0';
	
	signal bitvectord1319d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1319d : std_logic := '0';
	signal matchd1319d : std_logic := '0';
	
	signal bitvectord1320d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1320d : std_logic := '0';
	signal matchd1320d : std_logic := '0';
	
	signal bitvectord1321d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1321d : std_logic := '0';
	signal matchd1321d : std_logic := '0';
	
	signal bitvectord1322d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1322d : std_logic := '0';
	signal matchd1322d : std_logic := '0';
	
	signal bitvectord1323d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1323d : std_logic := '0';
	signal matchd1323d : std_logic := '0';
	
	signal bitvectord1324d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1324d : std_logic := '0';
	signal matchd1324d : std_logic := '0';
	
	signal bitvectord1325d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1325d : std_logic := '0';
	signal matchd1325d : std_logic := '0';
	
	signal bitvectord1326d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1326d : std_logic := '0';
	signal matchd1326d : std_logic := '0';
	
	signal bitvectord1327d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1327d : std_logic := '0';
	signal matchd1327d : std_logic := '0';
	
	signal bitvectord1328d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1328d : std_logic := '0';
	signal matchd1328d : std_logic := '0';
	
	signal bitvectord1329d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1329d : std_logic := '0';
	signal matchd1329d : std_logic := '0';
	
	signal bitvectord1330d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1330d : std_logic := '0';
	signal matchd1330d : std_logic := '0';
	
	signal bitvectord1331d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1331d : std_logic := '1';
	signal matchd1331d : std_logic := '0';
	
	signal bitvectord1332d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1332d : std_logic := '0';
	signal matchd1332d : std_logic := '0';
	
	signal bitvectord1333d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1333d : std_logic := '0';
	signal matchd1333d : std_logic := '0';
	
	signal bitvectord1334d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1334d : std_logic := '0';
	signal matchd1334d : std_logic := '0';
	
	signal bitvectord1335d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1335d : std_logic := '0';
	signal matchd1335d : std_logic := '0';
	
	signal bitvectord1336d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1336d : std_logic := '0';
	signal matchd1336d : std_logic := '0';
	
	signal bitvectord1337d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1337d : std_logic := '0';
	signal matchd1337d : std_logic := '0';
	
	signal bitvectord1338d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1338d : std_logic := '0';
	signal matchd1338d : std_logic := '0';
	
	signal bitvectord1339d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1339d : std_logic := '0';
	signal matchd1339d : std_logic := '0';
	
	signal bitvectord1340d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1340d : std_logic := '0';
	signal matchd1340d : std_logic := '0';
	
	signal bitvectord1341d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1341d : std_logic := '0';
	signal matchd1341d : std_logic := '0';
	
	signal bitvectord1342d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1342d : std_logic := '0';
	signal matchd1342d : std_logic := '0';
	
	signal bitvectord1343d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1343d : std_logic := '0';
	signal matchd1343d : std_logic := '0';
	
	signal bitvectord1344d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1344d : std_logic := '0';
	signal matchd1344d : std_logic := '0';
	
	signal bitvectord1345d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1345d : std_logic := '0';
	signal matchd1345d : std_logic := '0';
	
	signal bitvectord1346d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1346d : std_logic := '0';
	signal matchd1346d : std_logic := '0';
	
	signal bitvectord1347d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1347d : std_logic := '1';
	signal matchd1347d : std_logic := '0';
	
	signal bitvectord1348d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1348d : std_logic := '0';
	signal matchd1348d : std_logic := '0';
	
	signal bitvectord1349d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1349d : std_logic := '0';
	signal matchd1349d : std_logic := '0';
	
	signal bitvectord1350d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1350d : std_logic := '0';
	signal matchd1350d : std_logic := '0';
	
	signal bitvectord1351d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1351d : std_logic := '0';
	signal matchd1351d : std_logic := '0';
	
	signal bitvectord1352d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1352d : std_logic := '0';
	signal matchd1352d : std_logic := '0';
	
	signal bitvectord1353d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1353d : std_logic := '0';
	signal matchd1353d : std_logic := '0';
	
	signal bitvectord1354d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1354d : std_logic := '0';
	signal matchd1354d : std_logic := '0';
	
	signal bitvectord1355d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1355d : std_logic := '0';
	signal matchd1355d : std_logic := '0';
	
	signal bitvectord1356d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1356d : std_logic := '0';
	signal matchd1356d : std_logic := '0';
	
	signal bitvectord1357d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1357d : std_logic := '0';
	signal matchd1357d : std_logic := '0';
	
	signal bitvectord1358d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1358d : std_logic := '0';
	signal matchd1358d : std_logic := '0';
	
	signal bitvectord1359d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1359d : std_logic := '1';
	signal matchd1359d : std_logic := '0';
	
	signal bitvectord1360d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1360d : std_logic := '0';
	signal matchd1360d : std_logic := '0';
	
	signal bitvectord1361d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1361d : std_logic := '0';
	signal matchd1361d : std_logic := '0';
	
	signal bitvectord1362d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1362d : std_logic := '0';
	signal matchd1362d : std_logic := '0';
	
	signal bitvectord1363d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1363d : std_logic := '0';
	signal matchd1363d : std_logic := '0';
	
	signal bitvectord1364d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1364d : std_logic := '0';
	signal matchd1364d : std_logic := '0';
	
	signal bitvectord1365d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1365d : std_logic := '0';
	signal matchd1365d : std_logic := '0';
	
	signal bitvectord1366d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1366d : std_logic := '0';
	signal matchd1366d : std_logic := '0';
	
	signal bitvectord1367d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1367d : std_logic := '0';
	signal matchd1367d : std_logic := '0';
	
	signal bitvectord1368d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1368d : std_logic := '0';
	signal matchd1368d : std_logic := '0';
	
	signal bitvectord1369d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1369d : std_logic := '0';
	signal matchd1369d : std_logic := '0';
	
	signal bitvectord1370d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1370d : std_logic := '0';
	signal matchd1370d : std_logic := '0';
	
	signal bitvectord1371d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1371d : std_logic := '0';
	signal matchd1371d : std_logic := '0';
	
	signal bitvectord1372d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1372d : std_logic := '0';
	signal matchd1372d : std_logic := '0';
	
	signal bitvectord1373d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1373d : std_logic := '0';
	signal matchd1373d : std_logic := '0';
	
	signal bitvectord1374d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1374d : std_logic := '0';
	signal matchd1374d : std_logic := '0';
	
	signal bitvectord1375d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1375d : std_logic := '0';
	signal matchd1375d : std_logic := '0';
	
	signal bitvectord1376d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1376d : std_logic := '0';
	signal matchd1376d : std_logic := '0';
	
	signal bitvectord1377d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1377d : std_logic := '1';
	signal matchd1377d : std_logic := '0';
	
	signal bitvectord1378d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1378d : std_logic := '0';
	signal matchd1378d : std_logic := '0';
	
	signal bitvectord1379d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1379d : std_logic := '0';
	signal matchd1379d : std_logic := '0';
	
	signal bitvectord1380d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1380d : std_logic := '0';
	signal matchd1380d : std_logic := '0';
	
	signal bitvectord1381d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1381d : std_logic := '0';
	signal matchd1381d : std_logic := '0';
	
	signal bitvectord1382d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1382d : std_logic := '0';
	signal matchd1382d : std_logic := '0';
	
	signal bitvectord1383d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1383d : std_logic := '0';
	signal matchd1383d : std_logic := '0';
	
	signal bitvectord1384d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1384d : std_logic := '0';
	signal matchd1384d : std_logic := '0';
	
	signal bitvectord1385d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000";
	signal Enabled1385d : std_logic := '0';
	signal matchd1385d : std_logic := '0';
	
	signal bitvectord1386d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1386d : std_logic := '0';
	signal matchd1386d : std_logic := '0';
	
	signal bitvectord1387d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1387d : std_logic := '1';
	signal matchd1387d : std_logic := '0';
	
	signal bitvectord1388d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1388d : std_logic := '0';
	signal matchd1388d : std_logic := '0';
	
	signal bitvectord1389d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1389d : std_logic := '0';
	signal matchd1389d : std_logic := '0';
	
	signal bitvectord1390d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000";
	signal Enabled1390d : std_logic := '0';
	signal matchd1390d : std_logic := '0';
	
	signal bitvectord1391d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1391d : std_logic := '0';
	signal matchd1391d : std_logic := '0';
	
	signal bitvectord1392d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1392d : std_logic := '0';
	signal matchd1392d : std_logic := '0';
	
	signal bitvectord1393d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1393d : std_logic := '0';
	signal matchd1393d : std_logic := '0';
	
	signal bitvectord1394d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1394d : std_logic := '0';
	signal matchd1394d : std_logic := '0';
	
	signal bitvectord1395d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1395d : std_logic := '0';
	signal matchd1395d : std_logic := '0';
	
	signal bitvectord1396d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1396d : std_logic := '0';
	signal matchd1396d : std_logic := '0';
	
	signal bitvectord1397d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1397d : std_logic := '0';
	signal matchd1397d : std_logic := '0';
	
	signal bitvectord1398d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1398d : std_logic := '0';
	signal matchd1398d : std_logic := '0';
	
	signal bitvectord1399d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1399d : std_logic := '0';
	signal matchd1399d : std_logic := '0';
	
	signal bitvectord1400d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1400d : std_logic := '0';
	signal matchd1400d : std_logic := '0';
	
	signal bitvectord1401d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1401d : std_logic := '0';
	signal matchd1401d : std_logic := '0';
	
	signal bitvectord1402d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1402d : std_logic := '0';
	signal matchd1402d : std_logic := '0';
	
	signal bitvectord1403d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1403d : std_logic := '1';
	signal matchd1403d : std_logic := '0';
	
	signal bitvectord1404d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1404d : std_logic := '0';
	signal matchd1404d : std_logic := '0';
	
	signal bitvectord1405d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1405d : std_logic := '0';
	signal matchd1405d : std_logic := '0';
	
	signal bitvectord1406d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1406d : std_logic := '0';
	signal matchd1406d : std_logic := '0';
	
	signal bitvectord1407d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1407d : std_logic := '0';
	signal matchd1407d : std_logic := '0';
	
	signal bitvectord1408d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1408d : std_logic := '0';
	signal matchd1408d : std_logic := '0';
	
	signal bitvectord1409d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1409d : std_logic := '0';
	signal matchd1409d : std_logic := '0';
	
	signal bitvectord1410d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1410d : std_logic := '0';
	signal matchd1410d : std_logic := '0';
	
	signal bitvectord1411d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1411d : std_logic := '0';
	signal matchd1411d : std_logic := '0';
	
	signal bitvectord1412d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1412d : std_logic := '0';
	signal matchd1412d : std_logic := '0';
	
	signal bitvectord1413d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1413d : std_logic := '0';
	signal matchd1413d : std_logic := '0';
	
	signal bitvectord1414d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1414d : std_logic := '1';
	signal matchd1414d : std_logic := '0';
	
	signal bitvectord1415d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1415d : std_logic := '0';
	signal matchd1415d : std_logic := '0';
	
	signal bitvectord1416d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1416d : std_logic := '0';
	signal matchd1416d : std_logic := '0';
	
	signal bitvectord1417d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1417d : std_logic := '0';
	signal matchd1417d : std_logic := '0';
	
	signal bitvectord1418d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1418d : std_logic := '0';
	signal matchd1418d : std_logic := '0';
	
	signal bitvectord1419d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1419d : std_logic := '0';
	signal matchd1419d : std_logic := '0';
	
	signal bitvectord1420d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1420d : std_logic := '0';
	signal matchd1420d : std_logic := '0';
	
	signal bitvectord1421d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1421d : std_logic := '0';
	signal matchd1421d : std_logic := '0';
	
	signal bitvectord1422d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1422d : std_logic := '0';
	signal matchd1422d : std_logic := '0';
	
	signal bitvectord1423d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1423d : std_logic := '0';
	signal matchd1423d : std_logic := '0';
	
	signal bitvectord1424d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1424d : std_logic := '0';
	signal matchd1424d : std_logic := '0';
	
	signal bitvectord1425d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1425d : std_logic := '0';
	signal matchd1425d : std_logic := '0';
	
	signal bitvectord1426d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1426d : std_logic := '0';
	signal matchd1426d : std_logic := '0';
	
	signal bitvectord1427d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1427d : std_logic := '0';
	signal matchd1427d : std_logic := '0';
	
	signal bitvectord1428d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1428d : std_logic := '0';
	signal matchd1428d : std_logic := '0';
	
	signal bitvectord1429d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1429d : std_logic := '0';
	signal matchd1429d : std_logic := '0';
	
	signal bitvectord1430d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1430d : std_logic := '1';
	signal matchd1430d : std_logic := '0';
	
	signal bitvectord1431d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1431d : std_logic := '0';
	signal matchd1431d : std_logic := '0';
	
	signal bitvectord1432d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1432d : std_logic := '0';
	signal matchd1432d : std_logic := '0';
	
	signal bitvectord1433d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1433d : std_logic := '0';
	signal matchd1433d : std_logic := '0';
	
	signal bitvectord1434d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1434d : std_logic := '0';
	signal matchd1434d : std_logic := '0';
	
	signal bitvectord1435d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1435d : std_logic := '0';
	signal matchd1435d : std_logic := '0';
	
	signal bitvectord1436d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1436d : std_logic := '0';
	signal matchd1436d : std_logic := '0';
	
	signal bitvectord1437d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1437d : std_logic := '0';
	signal matchd1437d : std_logic := '0';
	
	signal bitvectord1438d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1438d : std_logic := '0';
	signal matchd1438d : std_logic := '0';
	
	signal bitvectord1439d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1439d : std_logic := '0';
	signal matchd1439d : std_logic := '0';
	
	signal bitvectord1440d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1440d : std_logic := '0';
	signal matchd1440d : std_logic := '0';
	
	signal bitvectord1441d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1441d : std_logic := '0';
	signal matchd1441d : std_logic := '0';
	
	signal bitvectord1442d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1442d : std_logic := '0';
	signal matchd1442d : std_logic := '0';
	
	signal bitvectord1443d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1443d : std_logic := '1';
	signal matchd1443d : std_logic := '0';
	
	signal bitvectord1444d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1444d : std_logic := '0';
	signal matchd1444d : std_logic := '0';
	
	signal bitvectord1445d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1445d : std_logic := '0';
	signal matchd1445d : std_logic := '0';
	
	signal bitvectord1446d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1446d : std_logic := '0';
	signal matchd1446d : std_logic := '0';
	
	signal bitvectord1447d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1447d : std_logic := '0';
	signal matchd1447d : std_logic := '0';
	
	signal bitvectord1448d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1448d : std_logic := '0';
	signal matchd1448d : std_logic := '0';
	
	signal bitvectord1449d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1449d : std_logic := '0';
	signal matchd1449d : std_logic := '0';
	
	signal bitvectord1450d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1450d : std_logic := '0';
	signal matchd1450d : std_logic := '0';
	
	signal bitvectord1451d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1451d : std_logic := '0';
	signal matchd1451d : std_logic := '0';
	
	signal bitvectord1452d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1452d : std_logic := '0';
	signal matchd1452d : std_logic := '0';
	
	signal bitvectord1453d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1453d : std_logic := '0';
	signal matchd1453d : std_logic := '0';
	
	signal bitvectord1454d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1454d : std_logic := '0';
	signal matchd1454d : std_logic := '0';
	
	signal bitvectord1455d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1455d : std_logic := '1';
	signal matchd1455d : std_logic := '0';
	
	signal bitvectord1456d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1456d : std_logic := '0';
	signal matchd1456d : std_logic := '0';
	
	signal bitvectord1457d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1457d : std_logic := '0';
	signal matchd1457d : std_logic := '0';
	
	signal bitvectord1458d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1458d : std_logic := '0';
	signal matchd1458d : std_logic := '0';
	
	signal bitvectord1459d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1459d : std_logic := '0';
	signal matchd1459d : std_logic := '0';
	
	signal bitvectord1460d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1460d : std_logic := '0';
	signal matchd1460d : std_logic := '0';
	
	signal bitvectord1461d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000";
	signal Enabled1461d : std_logic := '0';
	signal matchd1461d : std_logic := '0';
	
	signal bitvectord1462d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1462d : std_logic := '0';
	signal matchd1462d : std_logic := '0';
	
	signal bitvectord1463d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1463d : std_logic := '0';
	signal matchd1463d : std_logic := '0';
	
	signal bitvectord1464d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1464d : std_logic := '0';
	signal matchd1464d : std_logic := '0';
	
	signal bitvectord1465d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1465d : std_logic := '0';
	signal matchd1465d : std_logic := '0';
	
	signal bitvectord1466d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1466d : std_logic := '0';
	signal matchd1466d : std_logic := '0';
	
	signal bitvectord1467d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1467d : std_logic := '0';
	signal matchd1467d : std_logic := '0';
	
	signal bitvectord1468d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1468d : std_logic := '1';
	signal matchd1468d : std_logic := '0';
	
	signal bitvectord1469d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1469d : std_logic := '0';
	signal matchd1469d : std_logic := '0';
	
	signal bitvectord1470d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1470d : std_logic := '0';
	signal matchd1470d : std_logic := '0';
	
	signal bitvectord1471d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1471d : std_logic := '0';
	signal matchd1471d : std_logic := '0';
	
	signal bitvectord1472d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1472d : std_logic := '0';
	signal matchd1472d : std_logic := '0';
	
	signal bitvectord1473d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1473d : std_logic := '0';
	signal matchd1473d : std_logic := '0';
	
	signal bitvectord1474d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1474d : std_logic := '0';
	signal matchd1474d : std_logic := '0';
	
	signal bitvectord1475d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1475d : std_logic := '0';
	signal matchd1475d : std_logic := '0';
	
	signal bitvectord1476d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1476d : std_logic := '0';
	signal matchd1476d : std_logic := '0';
	
	signal bitvectord1477d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1477d : std_logic := '0';
	signal matchd1477d : std_logic := '0';
	
	signal bitvectord1478d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1478d : std_logic := '0';
	signal matchd1478d : std_logic := '0';
	
	signal bitvectord1479d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1479d : std_logic := '0';
	signal matchd1479d : std_logic := '0';
	
	signal bitvectord1480d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1480d : std_logic := '1';
	signal matchd1480d : std_logic := '0';
	
	signal bitvectord1481d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1481d : std_logic := '0';
	signal matchd1481d : std_logic := '0';
	
	signal bitvectord1482d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1482d : std_logic := '0';
	signal matchd1482d : std_logic := '0';
	
	signal bitvectord1483d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1483d : std_logic := '0';
	signal matchd1483d : std_logic := '0';
	
	signal bitvectord1484d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1484d : std_logic := '0';
	signal matchd1484d : std_logic := '0';
	
	signal bitvectord1485d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1485d : std_logic := '0';
	signal matchd1485d : std_logic := '0';
	
	signal bitvectord1486d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000";
	signal Enabled1486d : std_logic := '0';
	signal matchd1486d : std_logic := '0';
	
	signal bitvectord1487d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1487d : std_logic := '0';
	signal matchd1487d : std_logic := '0';
	
	signal bitvectord1488d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1488d : std_logic := '0';
	signal matchd1488d : std_logic := '0';
	
	signal bitvectord1489d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1489d : std_logic := '0';
	signal matchd1489d : std_logic := '0';
	
	signal bitvectord1490d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1490d : std_logic := '0';
	signal matchd1490d : std_logic := '0';
	
	signal bitvectord1491d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1491d : std_logic := '0';
	signal matchd1491d : std_logic := '0';
	
	signal bitvectord1492d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1492d : std_logic := '0';
	signal matchd1492d : std_logic := '0';
	
	signal bitvectord1493d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1493d : std_logic := '1';
	signal matchd1493d : std_logic := '0';
	
	signal bitvectord1494d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1494d : std_logic := '0';
	signal matchd1494d : std_logic := '0';
	
	signal bitvectord1495d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1495d : std_logic := '0';
	signal matchd1495d : std_logic := '0';
	
	signal bitvectord1496d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1496d : std_logic := '0';
	signal matchd1496d : std_logic := '0';
	
	signal bitvectord1497d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1497d : std_logic := '0';
	signal matchd1497d : std_logic := '0';
	
	signal bitvectord1498d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1498d : std_logic := '0';
	signal matchd1498d : std_logic := '0';
	
	signal bitvectord1499d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1499d : std_logic := '0';
	signal matchd1499d : std_logic := '0';
	
	signal bitvectord1500d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1500d : std_logic := '0';
	signal matchd1500d : std_logic := '0';
	
	signal bitvectord1501d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1501d : std_logic := '0';
	signal matchd1501d : std_logic := '0';
	
	signal bitvectord1502d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1502d : std_logic := '0';
	signal matchd1502d : std_logic := '0';
	
	signal bitvectord1503d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1503d : std_logic := '0';
	signal matchd1503d : std_logic := '0';
	
	signal bitvectord1504d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1504d : std_logic := '0';
	signal matchd1504d : std_logic := '0';
	
	signal bitvectord1505d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1505d : std_logic := '0';
	signal matchd1505d : std_logic := '0';
	
	signal bitvectord1506d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1506d : std_logic := '0';
	signal matchd1506d : std_logic := '0';
	
	signal bitvectord1507d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1507d : std_logic := '0';
	signal matchd1507d : std_logic := '0';
	
	signal bitvectord1508d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1508d : std_logic := '0';
	signal matchd1508d : std_logic := '0';
	
	signal bitvectord1509d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1509d : std_logic := '0';
	signal matchd1509d : std_logic := '0';
	
	signal bitvectord1510d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1510d : std_logic := '1';
	signal matchd1510d : std_logic := '0';
	
	signal bitvectord1511d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1511d : std_logic := '0';
	signal matchd1511d : std_logic := '0';
	
	signal bitvectord1512d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1512d : std_logic := '0';
	signal matchd1512d : std_logic := '0';
	
	signal bitvectord1513d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1513d : std_logic := '0';
	signal matchd1513d : std_logic := '0';
	
	signal bitvectord1514d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1514d : std_logic := '0';
	signal matchd1514d : std_logic := '0';
	
	signal bitvectord1515d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1515d : std_logic := '0';
	signal matchd1515d : std_logic := '0';
	
	signal bitvectord1516d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1516d : std_logic := '0';
	signal matchd1516d : std_logic := '0';
	
	signal bitvectord1517d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1517d : std_logic := '0';
	signal matchd1517d : std_logic := '0';
	
	signal bitvectord1518d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1518d : std_logic := '0';
	signal matchd1518d : std_logic := '0';
	
	signal bitvectord1519d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1519d : std_logic := '0';
	signal matchd1519d : std_logic := '0';
	
	signal bitvectord1520d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1520d : std_logic := '0';
	signal matchd1520d : std_logic := '0';
	
	signal bitvectord1521d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1521d : std_logic := '0';
	signal matchd1521d : std_logic := '0';
	
	signal bitvectord1522d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1522d : std_logic := '0';
	signal matchd1522d : std_logic := '0';
	
	signal bitvectord1523d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1523d : std_logic := '0';
	signal matchd1523d : std_logic := '0';
	
	signal bitvectord1524d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1524d : std_logic := '0';
	signal matchd1524d : std_logic := '0';
	
	signal bitvectord1525d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1525d : std_logic := '0';
	signal matchd1525d : std_logic := '0';
	
	signal bitvectord1526d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1526d : std_logic := '0';
	signal matchd1526d : std_logic := '0';
	
	signal bitvectord1527d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1527d : std_logic := '1';
	signal matchd1527d : std_logic := '0';
	
	signal bitvectord1528d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1528d : std_logic := '0';
	signal matchd1528d : std_logic := '0';
	
	signal bitvectord1529d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1529d : std_logic := '0';
	signal matchd1529d : std_logic := '0';
	
	signal bitvectord1530d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1530d : std_logic := '0';
	signal matchd1530d : std_logic := '0';
	
	signal bitvectord1531d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1531d : std_logic := '0';
	signal matchd1531d : std_logic := '0';
	
	signal bitvectord1532d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1532d : std_logic := '0';
	signal matchd1532d : std_logic := '0';
	
	signal bitvectord1533d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1533d : std_logic := '0';
	signal matchd1533d : std_logic := '0';
	
	signal bitvectord1534d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1534d : std_logic := '0';
	signal matchd1534d : std_logic := '0';
	
	signal bitvectord1535d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000";
	signal Enabled1535d : std_logic := '0';
	signal matchd1535d : std_logic := '0';
	
	signal bitvectord1536d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1536d : std_logic := '0';
	signal matchd1536d : std_logic := '0';
	
	signal bitvectord1537d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1537d : std_logic := '0';
	signal matchd1537d : std_logic := '0';
	
	signal bitvectord1538d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1538d : std_logic := '0';
	signal matchd1538d : std_logic := '0';
	
	signal bitvectord1539d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1539d : std_logic := '0';
	signal matchd1539d : std_logic := '0';
	
	signal bitvectord1540d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1540d : std_logic := '0';
	signal matchd1540d : std_logic := '0';
	
	signal bitvectord1541d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1541d : std_logic := '0';
	signal matchd1541d : std_logic := '0';
	
	signal bitvectord1542d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1542d : std_logic := '1';
	signal matchd1542d : std_logic := '0';
	
	signal bitvectord1543d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1543d : std_logic := '0';
	signal matchd1543d : std_logic := '0';
	
	signal bitvectord1544d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1544d : std_logic := '0';
	signal matchd1544d : std_logic := '0';
	
	signal bitvectord1545d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1545d : std_logic := '0';
	signal matchd1545d : std_logic := '0';
	
	signal bitvectord1546d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1546d : std_logic := '0';
	signal matchd1546d : std_logic := '0';
	
	signal bitvectord1547d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1547d : std_logic := '0';
	signal matchd1547d : std_logic := '0';
	
	signal bitvectord1548d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled1548d : std_logic := '0';
	signal matchd1548d : std_logic := '0';
	
	signal bitvectord1549d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1549d : std_logic := '0';
	signal matchd1549d : std_logic := '0';
	
	signal bitvectord1550d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1550d : std_logic := '0';
	signal matchd1550d : std_logic := '0';
	
	signal bitvectord1551d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1551d : std_logic := '0';
	signal matchd1551d : std_logic := '0';
	
	signal bitvectord1552d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1552d : std_logic := '0';
	signal matchd1552d : std_logic := '0';
	
	signal bitvectord1553d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1553d : std_logic := '0';
	signal matchd1553d : std_logic := '0';
	
	signal bitvectord1554d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1554d : std_logic := '0';
	signal matchd1554d : std_logic := '0';
	
	signal bitvectord1555d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1555d : std_logic := '0';
	signal matchd1555d : std_logic := '0';
	
	signal bitvectord1556d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1556d : std_logic := '1';
	signal matchd1556d : std_logic := '0';
	
	signal bitvectord1557d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1557d : std_logic := '0';
	signal matchd1557d : std_logic := '0';
	
	signal bitvectord1558d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1558d : std_logic := '0';
	signal matchd1558d : std_logic := '0';
	
	signal bitvectord1559d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1559d : std_logic := '0';
	signal matchd1559d : std_logic := '0';
	
	signal bitvectord1560d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1560d : std_logic := '0';
	signal matchd1560d : std_logic := '0';
	
	signal bitvectord1561d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1561d : std_logic := '0';
	signal matchd1561d : std_logic := '0';
	
	signal bitvectord1562d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1562d : std_logic := '0';
	signal matchd1562d : std_logic := '0';
	
	signal bitvectord1563d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1563d : std_logic := '0';
	signal matchd1563d : std_logic := '0';
	
	signal bitvectord1564d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1564d : std_logic := '0';
	signal matchd1564d : std_logic := '0';
	
	signal bitvectord1565d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1565d : std_logic := '0';
	signal matchd1565d : std_logic := '0';
	
	signal bitvectord1566d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1566d : std_logic := '0';
	signal matchd1566d : std_logic := '0';
	
	signal bitvectord1567d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1567d : std_logic := '0';
	signal matchd1567d : std_logic := '0';
	
	signal bitvectord1568d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1568d : std_logic := '0';
	signal matchd1568d : std_logic := '0';
	
	signal bitvectord1569d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1569d : std_logic := '0';
	signal matchd1569d : std_logic := '0';
	
	signal bitvectord1570d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1570d : std_logic := '0';
	signal matchd1570d : std_logic := '0';
	
	signal bitvectord1571d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1571d : std_logic := '0';
	signal matchd1571d : std_logic := '0';
	
	signal bitvectord1572d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1572d : std_logic := '0';
	signal matchd1572d : std_logic := '0';
	
	signal bitvectord1573d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1573d : std_logic := '1';
	signal matchd1573d : std_logic := '0';
	
	signal bitvectord1574d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1574d : std_logic := '0';
	signal matchd1574d : std_logic := '0';
	
	signal bitvectord1575d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1575d : std_logic := '0';
	signal matchd1575d : std_logic := '0';
	
	signal bitvectord1576d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1576d : std_logic := '0';
	signal matchd1576d : std_logic := '0';
	
	signal bitvectord1577d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1577d : std_logic := '0';
	signal matchd1577d : std_logic := '0';
	
	signal bitvectord1578d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1578d : std_logic := '0';
	signal matchd1578d : std_logic := '0';
	
	signal bitvectord1579d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1579d : std_logic := '0';
	signal matchd1579d : std_logic := '0';
	
	signal bitvectord1580d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1580d : std_logic := '0';
	signal matchd1580d : std_logic := '0';
	
	signal bitvectord1581d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1581d : std_logic := '0';
	signal matchd1581d : std_logic := '0';
	
	signal bitvectord1582d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1582d : std_logic := '0';
	signal matchd1582d : std_logic := '0';
	
	signal bitvectord1583d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1583d : std_logic := '0';
	signal matchd1583d : std_logic := '0';
	
	signal bitvectord1584d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1584d : std_logic := '0';
	signal matchd1584d : std_logic := '0';
	
	signal bitvectord1585d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1585d : std_logic := '1';
	signal matchd1585d : std_logic := '0';
	
	signal bitvectord1586d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1586d : std_logic := '0';
	signal matchd1586d : std_logic := '0';
	
	signal bitvectord1587d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1587d : std_logic := '0';
	signal matchd1587d : std_logic := '0';
	
	signal bitvectord1588d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1588d : std_logic := '0';
	signal matchd1588d : std_logic := '0';
	
	signal bitvectord1589d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1589d : std_logic := '0';
	signal matchd1589d : std_logic := '0';
	
	signal bitvectord1590d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1590d : std_logic := '0';
	signal matchd1590d : std_logic := '0';
	
	signal bitvectord1591d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1591d : std_logic := '0';
	signal matchd1591d : std_logic := '0';
	
	signal bitvectord1592d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1592d : std_logic := '0';
	signal matchd1592d : std_logic := '0';
	
	signal bitvectord1593d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1593d : std_logic := '0';
	signal matchd1593d : std_logic := '0';
	
	signal bitvectord1594d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1594d : std_logic := '0';
	signal matchd1594d : std_logic := '0';
	
	signal bitvectord1595d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1595d : std_logic := '0';
	signal matchd1595d : std_logic := '0';
	
	signal bitvectord1596d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1596d : std_logic := '0';
	signal matchd1596d : std_logic := '0';
	
	signal bitvectord1597d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1597d : std_logic := '0';
	signal matchd1597d : std_logic := '0';
	
	signal bitvectord1598d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1598d : std_logic := '0';
	signal matchd1598d : std_logic := '0';
	
	signal bitvectord1599d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1599d : std_logic := '1';
	signal matchd1599d : std_logic := '0';
	
	signal bitvectord1600d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1600d : std_logic := '0';
	signal matchd1600d : std_logic := '0';
	
	signal bitvectord1601d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1601d : std_logic := '0';
	signal matchd1601d : std_logic := '0';
	
	signal bitvectord1602d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1602d : std_logic := '0';
	signal matchd1602d : std_logic := '0';
	
	signal bitvectord1603d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1603d : std_logic := '0';
	signal matchd1603d : std_logic := '0';
	
	signal bitvectord1604d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1604d : std_logic := '0';
	signal matchd1604d : std_logic := '0';
	
	signal bitvectord1605d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1605d : std_logic := '0';
	signal matchd1605d : std_logic := '0';
	
	signal bitvectord1606d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1606d : std_logic := '0';
	signal matchd1606d : std_logic := '0';
	
	signal bitvectord1607d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1607d : std_logic := '0';
	signal matchd1607d : std_logic := '0';
	
	signal bitvectord1608d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1608d : std_logic := '0';
	signal matchd1608d : std_logic := '0';
	
	signal bitvectord1609d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1609d : std_logic := '0';
	signal matchd1609d : std_logic := '0';
	
	signal bitvectord1610d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1610d : std_logic := '1';
	signal matchd1610d : std_logic := '0';
	
	signal bitvectord1611d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1611d : std_logic := '0';
	signal matchd1611d : std_logic := '0';
	
	signal bitvectord1612d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1612d : std_logic := '0';
	signal matchd1612d : std_logic := '0';
	
	signal bitvectord1613d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1613d : std_logic := '0';
	signal matchd1613d : std_logic := '0';
	
	signal bitvectord1614d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1614d : std_logic := '0';
	signal matchd1614d : std_logic := '0';
	
	signal bitvectord1615d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1615d : std_logic := '0';
	signal matchd1615d : std_logic := '0';
	
	signal bitvectord1616d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1616d : std_logic := '0';
	signal matchd1616d : std_logic := '0';
	
	signal bitvectord1617d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1617d : std_logic := '0';
	signal matchd1617d : std_logic := '0';
	
	signal bitvectord1618d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1618d : std_logic := '0';
	signal matchd1618d : std_logic := '0';
	
	signal bitvectord1619d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1619d : std_logic := '0';
	signal matchd1619d : std_logic := '0';
	
	signal bitvectord1620d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1620d : std_logic := '0';
	signal matchd1620d : std_logic := '0';
	
	signal bitvectord1621d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1621d : std_logic := '0';
	signal matchd1621d : std_logic := '0';
	
	signal bitvectord1622d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1622d : std_logic := '1';
	signal matchd1622d : std_logic := '0';
	
	signal bitvectord1623d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1623d : std_logic := '0';
	signal matchd1623d : std_logic := '0';
	
	signal bitvectord1624d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1624d : std_logic := '0';
	signal matchd1624d : std_logic := '0';
	
	signal bitvectord1625d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1625d : std_logic := '0';
	signal matchd1625d : std_logic := '0';
	
	signal bitvectord1626d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1626d : std_logic := '0';
	signal matchd1626d : std_logic := '0';
	
	signal bitvectord1627d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1627d : std_logic := '0';
	signal matchd1627d : std_logic := '0';
	
	signal bitvectord1628d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1628d : std_logic := '0';
	signal matchd1628d : std_logic := '0';
	
	signal bitvectord1629d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1629d : std_logic := '0';
	signal matchd1629d : std_logic := '0';
	
	signal bitvectord1630d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1630d : std_logic := '0';
	signal matchd1630d : std_logic := '0';
	
	signal bitvectord1631d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1631d : std_logic := '1';
	signal matchd1631d : std_logic := '0';
	
	signal bitvectord1632d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1632d : std_logic := '0';
	signal matchd1632d : std_logic := '0';
	
	signal bitvectord1633d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1633d : std_logic := '0';
	signal matchd1633d : std_logic := '0';
	
	signal bitvectord1634d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1634d : std_logic := '0';
	signal matchd1634d : std_logic := '0';
	
	signal bitvectord1635d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1635d : std_logic := '0';
	signal matchd1635d : std_logic := '0';
	
	signal bitvectord1636d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1636d : std_logic := '0';
	signal matchd1636d : std_logic := '0';
	
	signal bitvectord1637d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1637d : std_logic := '0';
	signal matchd1637d : std_logic := '0';
	
	signal bitvectord1638d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1638d : std_logic := '0';
	signal matchd1638d : std_logic := '0';
	
	signal bitvectord1639d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1639d : std_logic := '0';
	signal matchd1639d : std_logic := '0';
	
	signal bitvectord1640d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1640d : std_logic := '0';
	signal matchd1640d : std_logic := '0';
	
	signal bitvectord1641d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1641d : std_logic := '0';
	signal matchd1641d : std_logic := '0';
	
	signal bitvectord1642d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1642d : std_logic := '0';
	signal matchd1642d : std_logic := '0';
	
	signal bitvectord1643d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1643d : std_logic := '1';
	signal matchd1643d : std_logic := '0';
	
	signal bitvectord1644d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1644d : std_logic := '0';
	signal matchd1644d : std_logic := '0';
	
	signal bitvectord1645d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1645d : std_logic := '0';
	signal matchd1645d : std_logic := '0';
	
	signal bitvectord1646d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1646d : std_logic := '0';
	signal matchd1646d : std_logic := '0';
	
	signal bitvectord1647d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1647d : std_logic := '0';
	signal matchd1647d : std_logic := '0';
	
	signal bitvectord1648d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1648d : std_logic := '0';
	signal matchd1648d : std_logic := '0';
	
	signal bitvectord1649d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1649d : std_logic := '0';
	signal matchd1649d : std_logic := '0';
	
	signal bitvectord1650d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1650d : std_logic := '0';
	signal matchd1650d : std_logic := '0';
	
	signal bitvectord1651d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1651d : std_logic := '0';
	signal matchd1651d : std_logic := '0';
	
	signal bitvectord1652d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1652d : std_logic := '0';
	signal matchd1652d : std_logic := '0';
	
	signal bitvectord1653d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1653d : std_logic := '0';
	signal matchd1653d : std_logic := '0';
	
	signal bitvectord1654d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1654d : std_logic := '1';
	signal matchd1654d : std_logic := '0';
	
	signal bitvectord1655d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1655d : std_logic := '0';
	signal matchd1655d : std_logic := '0';
	
	signal bitvectord1656d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1656d : std_logic := '0';
	signal matchd1656d : std_logic := '0';
	
	signal bitvectord1657d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1657d : std_logic := '0';
	signal matchd1657d : std_logic := '0';
	
	signal bitvectord1658d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1658d : std_logic := '0';
	signal matchd1658d : std_logic := '0';
	
	signal bitvectord1659d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1659d : std_logic := '0';
	signal matchd1659d : std_logic := '0';
	
	signal bitvectord1660d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1660d : std_logic := '0';
	signal matchd1660d : std_logic := '0';
	
	signal bitvectord1661d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1661d : std_logic := '0';
	signal matchd1661d : std_logic := '0';
	
	signal bitvectord1662d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1662d : std_logic := '0';
	signal matchd1662d : std_logic := '0';
	
	signal bitvectord1663d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1663d : std_logic := '0';
	signal matchd1663d : std_logic := '0';
	
	signal bitvectord1664d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1664d : std_logic := '0';
	signal matchd1664d : std_logic := '0';
	
	signal bitvectord1665d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1665d : std_logic := '0';
	signal matchd1665d : std_logic := '0';
	
	signal bitvectord1666d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1666d : std_logic := '0';
	signal matchd1666d : std_logic := '0';
	
	signal bitvectord1667d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1667d : std_logic := '0';
	signal matchd1667d : std_logic := '0';
	
	signal bitvectord1668d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1668d : std_logic := '0';
	signal matchd1668d : std_logic := '0';
	
	signal bitvectord1669d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1669d : std_logic := '0';
	signal matchd1669d : std_logic := '0';
	
	signal bitvectord1670d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1670d : std_logic := '0';
	signal matchd1670d : std_logic := '0';
	
	signal bitvectord1671d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111";
	signal Enabled1671d : std_logic := '0';
	signal matchd1671d : std_logic := '0';
	
	signal bitvectord1672d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1672d : std_logic := '0';
	signal matchd1672d : std_logic := '0';
	
	signal bitvectord1673d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1673d : std_logic := '1';
	signal matchd1673d : std_logic := '0';
	
	signal bitvectord1674d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1674d : std_logic := '0';
	signal matchd1674d : std_logic := '0';
	
	signal bitvectord1675d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1675d : std_logic := '0';
	signal matchd1675d : std_logic := '0';
	
	signal bitvectord1676d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1676d : std_logic := '0';
	signal matchd1676d : std_logic := '0';
	
	signal bitvectord1677d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1677d : std_logic := '0';
	signal matchd1677d : std_logic := '0';
	
	signal bitvectord1678d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1678d : std_logic := '0';
	signal matchd1678d : std_logic := '0';
	
	signal bitvectord1679d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1679d : std_logic := '0';
	signal matchd1679d : std_logic := '0';
	
	signal bitvectord1680d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1680d : std_logic := '0';
	signal matchd1680d : std_logic := '0';
	
	signal bitvectord1681d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1681d : std_logic := '0';
	signal matchd1681d : std_logic := '0';
	
	signal bitvectord1682d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1682d : std_logic := '0';
	signal matchd1682d : std_logic := '0';
	
	signal bitvectord1683d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1683d : std_logic := '0';
	signal matchd1683d : std_logic := '0';
	
	signal bitvectord1684d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1684d : std_logic := '0';
	signal matchd1684d : std_logic := '0';
	
	signal bitvectord1685d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1685d : std_logic := '0';
	signal matchd1685d : std_logic := '0';
	
	signal bitvectord1686d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1686d : std_logic := '0';
	signal matchd1686d : std_logic := '0';
	
	signal bitvectord1687d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1687d : std_logic := '0';
	signal matchd1687d : std_logic := '0';
	
	signal bitvectord1688d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1688d : std_logic := '0';
	signal matchd1688d : std_logic := '0';
	
	signal bitvectord1689d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1689d : std_logic := '0';
	signal matchd1689d : std_logic := '0';
	
	signal bitvectord1690d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1690d : std_logic := '0';
	signal matchd1690d : std_logic := '0';
	
	signal bitvectord1691d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1691d : std_logic := '1';
	signal matchd1691d : std_logic := '0';
	
	signal bitvectord1692d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1692d : std_logic := '0';
	signal matchd1692d : std_logic := '0';
	
	signal bitvectord1693d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1693d : std_logic := '0';
	signal matchd1693d : std_logic := '0';
	
	signal bitvectord1694d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1694d : std_logic := '0';
	signal matchd1694d : std_logic := '0';
	
	signal bitvectord1695d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1695d : std_logic := '0';
	signal matchd1695d : std_logic := '0';
	
	signal bitvectord1696d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1696d : std_logic := '0';
	signal matchd1696d : std_logic := '0';
	
	signal bitvectord1697d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1697d : std_logic := '0';
	signal matchd1697d : std_logic := '0';
	
	signal bitvectord1698d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1698d : std_logic := '0';
	signal matchd1698d : std_logic := '0';
	
	signal bitvectord1699d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1699d : std_logic := '0';
	signal matchd1699d : std_logic := '0';
	
	signal bitvectord1700d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1700d : std_logic := '0';
	signal matchd1700d : std_logic := '0';
	
	signal bitvectord1701d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1701d : std_logic := '0';
	signal matchd1701d : std_logic := '0';
	
	signal bitvectord1702d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1702d : std_logic := '1';
	signal matchd1702d : std_logic := '0';
	
	signal bitvectord1703d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1703d : std_logic := '0';
	signal matchd1703d : std_logic := '0';
	
	signal bitvectord1704d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1704d : std_logic := '0';
	signal matchd1704d : std_logic := '0';
	
	signal bitvectord1705d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1705d : std_logic := '0';
	signal matchd1705d : std_logic := '0';
	
	signal bitvectord1706d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1706d : std_logic := '0';
	signal matchd1706d : std_logic := '0';
	
	signal bitvectord1707d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1707d : std_logic := '0';
	signal matchd1707d : std_logic := '0';
	
	signal bitvectord1708d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1708d : std_logic := '0';
	signal matchd1708d : std_logic := '0';
	
	signal bitvectord1709d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1709d : std_logic := '0';
	signal matchd1709d : std_logic := '0';
	
	signal bitvectord1710d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1710d : std_logic := '0';
	signal matchd1710d : std_logic := '0';
	
	signal bitvectord1711d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1711d : std_logic := '0';
	signal matchd1711d : std_logic := '0';
	
	signal bitvectord1712d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1712d : std_logic := '0';
	signal matchd1712d : std_logic := '0';
	
	signal bitvectord1713d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1713d : std_logic := '0';
	signal matchd1713d : std_logic := '0';
	
	signal bitvectord1714d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1714d : std_logic := '0';
	signal matchd1714d : std_logic := '0';
	
	signal bitvectord1715d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111";
	signal Enabled1715d : std_logic := '0';
	signal matchd1715d : std_logic := '0';
	
	signal bitvectord1716d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1716d : std_logic := '0';
	signal matchd1716d : std_logic := '0';
	
	signal bitvectord1717d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1717d : std_logic := '1';
	signal matchd1717d : std_logic := '0';
	
	signal bitvectord1718d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1718d : std_logic := '0';
	signal matchd1718d : std_logic := '0';
	
	signal bitvectord1719d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1719d : std_logic := '0';
	signal matchd1719d : std_logic := '0';
	
	signal bitvectord1720d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1720d : std_logic := '0';
	signal matchd1720d : std_logic := '0';
	
	signal bitvectord1721d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1721d : std_logic := '0';
	signal matchd1721d : std_logic := '0';
	
	signal bitvectord1722d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1722d : std_logic := '0';
	signal matchd1722d : std_logic := '0';
	
	signal bitvectord1723d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1723d : std_logic := '0';
	signal matchd1723d : std_logic := '0';
	
	signal bitvectord1724d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1724d : std_logic := '0';
	signal matchd1724d : std_logic := '0';
	
	signal bitvectord1725d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1725d : std_logic := '0';
	signal matchd1725d : std_logic := '0';
	
	signal bitvectord1726d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1726d : std_logic := '0';
	signal matchd1726d : std_logic := '0';
	
	signal bitvectord1727d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1727d : std_logic := '0';
	signal matchd1727d : std_logic := '0';
	
	signal bitvectord1728d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1728d : std_logic := '0';
	signal matchd1728d : std_logic := '0';
	
	signal bitvectord1729d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1729d : std_logic := '1';
	signal matchd1729d : std_logic := '0';
	
	signal bitvectord1730d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1730d : std_logic := '0';
	signal matchd1730d : std_logic := '0';
	
	signal bitvectord1731d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1731d : std_logic := '0';
	signal matchd1731d : std_logic := '0';
	
	signal bitvectord1732d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled1732d : std_logic := '0';
	signal matchd1732d : std_logic := '0';
	
	signal bitvectord1733d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1733d : std_logic := '0';
	signal matchd1733d : std_logic := '0';
	
	signal bitvectord1734d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1734d : std_logic := '0';
	signal matchd1734d : std_logic := '0';
	
	signal bitvectord1735d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1735d : std_logic := '0';
	signal matchd1735d : std_logic := '0';
	
	signal bitvectord1736d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1736d : std_logic := '0';
	signal matchd1736d : std_logic := '0';
	
	signal bitvectord1737d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1737d : std_logic := '0';
	signal matchd1737d : std_logic := '0';
	
	signal bitvectord1738d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1738d : std_logic := '0';
	signal matchd1738d : std_logic := '0';
	
	signal bitvectord1739d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled1739d : std_logic := '0';
	signal matchd1739d : std_logic := '0';
	
	signal bitvectord1740d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1740d : std_logic := '0';
	signal matchd1740d : std_logic := '0';
	
	signal bitvectord1741d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1741d : std_logic := '0';
	signal matchd1741d : std_logic := '0';
	
	signal bitvectord1742d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1742d : std_logic := '0';
	signal matchd1742d : std_logic := '0';
	
	signal bitvectord1743d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1743d : std_logic := '0';
	signal matchd1743d : std_logic := '0';
	
	signal bitvectord1744d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1744d : std_logic := '0';
	signal matchd1744d : std_logic := '0';
	
	signal bitvectord1745d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1745d : std_logic := '0';
	signal matchd1745d : std_logic := '0';
	
	signal bitvectord1746d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1746d : std_logic := '1';
	signal matchd1746d : std_logic := '0';
	
	signal bitvectord1747d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1747d : std_logic := '0';
	signal matchd1747d : std_logic := '0';
	
	signal bitvectord1748d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1748d : std_logic := '0';
	signal matchd1748d : std_logic := '0';
	
	signal bitvectord1749d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1749d : std_logic := '0';
	signal matchd1749d : std_logic := '0';
	
	signal bitvectord1750d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1750d : std_logic := '0';
	signal matchd1750d : std_logic := '0';
	
	signal bitvectord1751d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1751d : std_logic := '0';
	signal matchd1751d : std_logic := '0';
	
	signal bitvectord1752d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled1752d : std_logic := '0';
	signal matchd1752d : std_logic := '0';
	
	signal bitvectord1753d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1753d : std_logic := '0';
	signal matchd1753d : std_logic := '0';
	
	signal bitvectord1754d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1754d : std_logic := '0';
	signal matchd1754d : std_logic := '0';
	
	signal bitvectord1755d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1755d : std_logic := '0';
	signal matchd1755d : std_logic := '0';
	
	signal bitvectord1756d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled1756d : std_logic := '0';
	signal matchd1756d : std_logic := '0';
	
	signal bitvectord1757d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1757d : std_logic := '0';
	signal matchd1757d : std_logic := '0';
	
	signal bitvectord1758d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1758d : std_logic := '0';
	signal matchd1758d : std_logic := '0';
	
	signal bitvectord1759d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1759d : std_logic := '0';
	signal matchd1759d : std_logic := '0';
	
	signal bitvectord1760d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1760d : std_logic := '0';
	signal matchd1760d : std_logic := '0';
	
	signal bitvectord1761d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1761d : std_logic := '0';
	signal matchd1761d : std_logic := '0';
	
	signal bitvectord1762d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1762d : std_logic := '0';
	signal matchd1762d : std_logic := '0';
	
	signal bitvectord1764d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1764d : std_logic := '1';
	signal matchd1764d : std_logic := '0';
	
	signal bitvectord1765d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1765d : std_logic := '0';
	signal matchd1765d : std_logic := '0';
	
	signal bitvectord1766d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1766d : std_logic := '0';
	signal matchd1766d : std_logic := '0';
	
	signal bitvectord1767d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1767d : std_logic := '0';
	signal matchd1767d : std_logic := '0';
	
	signal bitvectord1768d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1768d : std_logic := '0';
	signal matchd1768d : std_logic := '0';
	
	signal bitvectord1769d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1769d : std_logic := '0';
	signal matchd1769d : std_logic := '0';
	
	signal bitvectord1770d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1770d : std_logic := '0';
	signal matchd1770d : std_logic := '0';
	
	signal bitvectord1771d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1771d : std_logic := '0';
	signal matchd1771d : std_logic := '0';
	
	signal bitvectord1772d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1772d : std_logic := '0';
	signal matchd1772d : std_logic := '0';
	
	signal bitvectord1773d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1773d : std_logic := '0';
	signal matchd1773d : std_logic := '0';
	
	signal bitvectord1774d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1774d : std_logic := '0';
	signal matchd1774d : std_logic := '0';
	
	signal bitvectord1775d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1775d : std_logic := '1';
	signal matchd1775d : std_logic := '0';
	
	signal bitvectord1776d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1776d : std_logic := '0';
	signal matchd1776d : std_logic := '0';
	
	signal bitvectord1777d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1777d : std_logic := '0';
	signal matchd1777d : std_logic := '0';
	
	signal bitvectord1778d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1778d : std_logic := '0';
	signal matchd1778d : std_logic := '0';
	
	signal bitvectord1779d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1779d : std_logic := '0';
	signal matchd1779d : std_logic := '0';
	
	signal bitvectord1780d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1780d : std_logic := '0';
	signal matchd1780d : std_logic := '0';
	
	signal bitvectord1781d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1781d : std_logic := '0';
	signal matchd1781d : std_logic := '0';
	
	signal bitvectord1782d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1782d : std_logic := '0';
	signal matchd1782d : std_logic := '0';
	
	signal bitvectord1783d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1783d : std_logic := '0';
	signal matchd1783d : std_logic := '0';
	
	signal bitvectord1784d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1784d : std_logic := '0';
	signal matchd1784d : std_logic := '0';
	
	signal bitvectord1785d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1785d : std_logic := '0';
	signal matchd1785d : std_logic := '0';
	
	signal bitvectord1786d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1786d : std_logic := '0';
	signal matchd1786d : std_logic := '0';
	
	signal bitvectord1787d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1787d : std_logic := '0';
	signal matchd1787d : std_logic := '0';
	
	signal bitvectord1788d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1788d : std_logic := '0';
	signal matchd1788d : std_logic := '0';
	
	signal bitvectord1789d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1789d : std_logic := '0';
	signal matchd1789d : std_logic := '0';
	
	signal bitvectord1790d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1790d : std_logic := '0';
	signal matchd1790d : std_logic := '0';
	
	signal bitvectord1791d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1791d : std_logic := '0';
	signal matchd1791d : std_logic := '0';
	
	signal bitvectord1792d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1792d : std_logic := '0';
	signal matchd1792d : std_logic := '0';
	
	signal bitvectord1793d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1793d : std_logic := '0';
	signal matchd1793d : std_logic := '0';
	
	signal bitvectord1794d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1794d : std_logic := '0';
	signal matchd1794d : std_logic := '0';
	
	signal bitvectord1795d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1795d : std_logic := '0';
	signal matchd1795d : std_logic := '0';
	
	signal bitvectord1796d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1796d : std_logic := '0';
	signal matchd1796d : std_logic := '0';
	
	signal bitvectord1797d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1797d : std_logic := '1';
	signal matchd1797d : std_logic := '0';
	
	signal bitvectord1798d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1798d : std_logic := '0';
	signal matchd1798d : std_logic := '0';
	
	signal bitvectord1799d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1799d : std_logic := '0';
	signal matchd1799d : std_logic := '0';
	
	signal bitvectord1800d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1800d : std_logic := '0';
	signal matchd1800d : std_logic := '0';
	
	signal bitvectord1801d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1801d : std_logic := '0';
	signal matchd1801d : std_logic := '0';
	
	signal bitvectord1802d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1802d : std_logic := '0';
	signal matchd1802d : std_logic := '0';
	
	signal bitvectord1803d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1803d : std_logic := '0';
	signal matchd1803d : std_logic := '0';
	
	signal bitvectord1804d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1804d : std_logic := '0';
	signal matchd1804d : std_logic := '0';
	
	signal bitvectord1805d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111";
	signal Enabled1805d : std_logic := '0';
	signal matchd1805d : std_logic := '0';
	
	signal bitvectord1806d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1806d : std_logic := '0';
	signal matchd1806d : std_logic := '0';
	
	signal bitvectord1807d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1807d : std_logic := '0';
	signal matchd1807d : std_logic := '0';
	
	signal bitvectord1808d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1808d : std_logic := '0';
	signal matchd1808d : std_logic := '0';
	
	signal bitvectord1809d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled1809d : std_logic := '0';
	signal matchd1809d : std_logic := '0';
	
	signal bitvectord1810d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1810d : std_logic := '0';
	signal matchd1810d : std_logic := '0';
	
	signal bitvectord1811d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1811d : std_logic := '0';
	signal matchd1811d : std_logic := '0';
	
	signal bitvectord1812d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1812d : std_logic := '0';
	signal matchd1812d : std_logic := '0';
	
	signal bitvectord1813d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled1813d : std_logic := '0';
	signal matchd1813d : std_logic := '0';
	
	signal bitvectord1814d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1814d : std_logic := '0';
	signal matchd1814d : std_logic := '0';
	
	signal bitvectord1815d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1815d : std_logic := '1';
	signal matchd1815d : std_logic := '0';
	
	signal bitvectord1816d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1816d : std_logic := '0';
	signal matchd1816d : std_logic := '0';
	
	signal bitvectord1817d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1817d : std_logic := '0';
	signal matchd1817d : std_logic := '0';
	
	signal bitvectord1818d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1818d : std_logic := '0';
	signal matchd1818d : std_logic := '0';
	
	signal bitvectord1819d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1819d : std_logic := '0';
	signal matchd1819d : std_logic := '0';
	
	signal bitvectord1820d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1820d : std_logic := '0';
	signal matchd1820d : std_logic := '0';
	
	signal bitvectord1821d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1821d : std_logic := '0';
	signal matchd1821d : std_logic := '0';
	
	signal bitvectord1822d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1822d : std_logic := '0';
	signal matchd1822d : std_logic := '0';
	
	signal bitvectord1823d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled1823d : std_logic := '0';
	signal matchd1823d : std_logic := '0';
	
	signal bitvectord1824d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1824d : std_logic := '0';
	signal matchd1824d : std_logic := '0';
	
	signal bitvectord1825d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1825d : std_logic := '0';
	signal matchd1825d : std_logic := '0';
	
	signal bitvectord1826d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1826d : std_logic := '0';
	signal matchd1826d : std_logic := '0';
	
	signal bitvectord1827d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111";
	signal Enabled1827d : std_logic := '0';
	signal matchd1827d : std_logic := '0';
	
	signal bitvectord1828d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1828d : std_logic := '0';
	signal matchd1828d : std_logic := '0';
	
	signal bitvectord1829d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1829d : std_logic := '0';
	signal matchd1829d : std_logic := '0';
	
	signal bitvectord1830d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1830d : std_logic := '0';
	signal matchd1830d : std_logic := '0';
	
	signal bitvectord1831d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled1831d : std_logic := '0';
	signal matchd1831d : std_logic := '0';
	
	signal bitvectord1832d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1832d : std_logic := '0';
	signal matchd1832d : std_logic := '0';
	
	signal bitvectord1833d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1833d : std_logic := '1';
	signal matchd1833d : std_logic := '0';
	
	signal bitvectord1834d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1834d : std_logic := '0';
	signal matchd1834d : std_logic := '0';
	
	signal bitvectord1835d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1835d : std_logic := '0';
	signal matchd1835d : std_logic := '0';
	
	signal bitvectord1836d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1836d : std_logic := '0';
	signal matchd1836d : std_logic := '0';
	
	signal bitvectord1837d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1837d : std_logic := '0';
	signal matchd1837d : std_logic := '0';
	
	signal bitvectord1838d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1838d : std_logic := '0';
	signal matchd1838d : std_logic := '0';
	
	signal bitvectord1839d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1839d : std_logic := '0';
	signal matchd1839d : std_logic := '0';
	
	signal bitvectord1840d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1840d : std_logic := '0';
	signal matchd1840d : std_logic := '0';
	
	signal bitvectord1841d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled1841d : std_logic := '0';
	signal matchd1841d : std_logic := '0';
	
	signal bitvectord1842d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1842d : std_logic := '0';
	signal matchd1842d : std_logic := '0';
	
	signal bitvectord1843d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1843d : std_logic := '0';
	signal matchd1843d : std_logic := '0';
	
	signal bitvectord1844d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1844d : std_logic := '0';
	signal matchd1844d : std_logic := '0';
	
	signal bitvectord1845d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled1845d : std_logic := '0';
	signal matchd1845d : std_logic := '0';
	
	signal bitvectord1846d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1846d : std_logic := '0';
	signal matchd1846d : std_logic := '0';
	
	signal bitvectord1847d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1847d : std_logic := '0';
	signal matchd1847d : std_logic := '0';
	
	signal bitvectord1848d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1848d : std_logic := '0';
	signal matchd1848d : std_logic := '0';
	
	signal bitvectord1849d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111";
	signal Enabled1849d : std_logic := '0';
	signal matchd1849d : std_logic := '0';
	
	signal bitvectord1850d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1850d : std_logic := '0';
	signal matchd1850d : std_logic := '0';
	
	signal bitvectord1852d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1852d : std_logic := '1';
	signal matchd1852d : std_logic := '0';
	
	signal bitvectord1853d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1853d : std_logic := '0';
	signal matchd1853d : std_logic := '0';
	
	signal bitvectord1854d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1854d : std_logic := '0';
	signal matchd1854d : std_logic := '0';
	
	signal bitvectord1855d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1855d : std_logic := '0';
	signal matchd1855d : std_logic := '0';
	
	signal bitvectord1856d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1856d : std_logic := '0';
	signal matchd1856d : std_logic := '0';
	
	signal bitvectord1857d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1857d : std_logic := '0';
	signal matchd1857d : std_logic := '0';
	
	signal bitvectord1858d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1858d : std_logic := '0';
	signal matchd1858d : std_logic := '0';
	
	signal bitvectord1859d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1859d : std_logic := '0';
	signal matchd1859d : std_logic := '0';
	
	signal bitvectord1860d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1860d : std_logic := '0';
	signal matchd1860d : std_logic := '0';
	
	signal bitvectord1861d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1861d : std_logic := '0';
	signal matchd1861d : std_logic := '0';
	
	signal bitvectord1862d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1862d : std_logic := '0';
	signal matchd1862d : std_logic := '0';
	
	signal bitvectord1863d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1863d : std_logic := '1';
	signal matchd1863d : std_logic := '0';
	
	signal bitvectord1864d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1864d : std_logic := '0';
	signal matchd1864d : std_logic := '0';
	
	signal bitvectord1865d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1865d : std_logic := '0';
	signal matchd1865d : std_logic := '0';
	
	signal bitvectord1866d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1866d : std_logic := '0';
	signal matchd1866d : std_logic := '0';
	
	signal bitvectord1867d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1867d : std_logic := '0';
	signal matchd1867d : std_logic := '0';
	
	signal bitvectord1868d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1868d : std_logic := '0';
	signal matchd1868d : std_logic := '0';
	
	signal bitvectord1869d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1869d : std_logic := '0';
	signal matchd1869d : std_logic := '0';
	
	signal bitvectord1870d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1870d : std_logic := '0';
	signal matchd1870d : std_logic := '0';
	
	signal bitvectord1871d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1871d : std_logic := '0';
	signal matchd1871d : std_logic := '0';
	
	signal bitvectord1872d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1872d : std_logic := '0';
	signal matchd1872d : std_logic := '0';
	
	signal bitvectord1873d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1873d : std_logic := '0';
	signal matchd1873d : std_logic := '0';
	
	signal bitvectord1874d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1874d : std_logic := '0';
	signal matchd1874d : std_logic := '0';
	
	signal bitvectord1875d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1875d : std_logic := '1';
	signal matchd1875d : std_logic := '0';
	
	signal bitvectord1876d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1876d : std_logic := '0';
	signal matchd1876d : std_logic := '0';
	
	signal bitvectord1877d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1877d : std_logic := '0';
	signal matchd1877d : std_logic := '0';
	
	signal bitvectord1878d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1878d : std_logic := '0';
	signal matchd1878d : std_logic := '0';
	
	signal bitvectord1879d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1879d : std_logic := '0';
	signal matchd1879d : std_logic := '0';
	
	signal bitvectord1880d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1880d : std_logic := '0';
	signal matchd1880d : std_logic := '0';
	
	signal bitvectord1881d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1881d : std_logic := '0';
	signal matchd1881d : std_logic := '0';
	
	signal bitvectord1882d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1882d : std_logic := '0';
	signal matchd1882d : std_logic := '0';
	
	signal bitvectord1883d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1883d : std_logic := '0';
	signal matchd1883d : std_logic := '0';
	
	signal bitvectord1884d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1884d : std_logic := '0';
	signal matchd1884d : std_logic := '0';
	
	signal bitvectord1885d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1885d : std_logic := '0';
	signal matchd1885d : std_logic := '0';
	
	signal bitvectord1886d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1886d : std_logic := '0';
	signal matchd1886d : std_logic := '0';
	
	signal bitvectord1887d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1887d : std_logic := '0';
	signal matchd1887d : std_logic := '0';
	
	signal bitvectord1888d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1888d : std_logic := '0';
	signal matchd1888d : std_logic := '0';
	
	signal bitvectord1889d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1889d : std_logic := '1';
	signal matchd1889d : std_logic := '0';
	
	signal bitvectord1890d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1890d : std_logic := '0';
	signal matchd1890d : std_logic := '0';
	
	signal bitvectord1891d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1891d : std_logic := '0';
	signal matchd1891d : std_logic := '0';
	
	signal bitvectord1892d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1892d : std_logic := '0';
	signal matchd1892d : std_logic := '0';
	
	signal bitvectord1893d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1893d : std_logic := '0';
	signal matchd1893d : std_logic := '0';
	
	signal bitvectord1894d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1894d : std_logic := '0';
	signal matchd1894d : std_logic := '0';
	
	signal bitvectord1895d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1895d : std_logic := '0';
	signal matchd1895d : std_logic := '0';
	
	signal bitvectord1896d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1896d : std_logic := '0';
	signal matchd1896d : std_logic := '0';
	
	signal bitvectord1897d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1897d : std_logic := '0';
	signal matchd1897d : std_logic := '0';
	
	signal bitvectord1898d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1898d : std_logic := '0';
	signal matchd1898d : std_logic := '0';
	
	signal bitvectord1899d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1899d : std_logic := '0';
	signal matchd1899d : std_logic := '0';
	
	signal bitvectord1900d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1900d : std_logic := '0';
	signal matchd1900d : std_logic := '0';
	
	signal bitvectord1901d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1901d : std_logic := '0';
	signal matchd1901d : std_logic := '0';
	
	signal bitvectord1902d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1902d : std_logic := '0';
	signal matchd1902d : std_logic := '0';
	
	signal bitvectord1903d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1903d : std_logic := '0';
	signal matchd1903d : std_logic := '0';
	
	signal bitvectord1904d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1904d : std_logic := '0';
	signal matchd1904d : std_logic := '0';
	
	signal bitvectord1905d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1905d : std_logic := '1';
	signal matchd1905d : std_logic := '0';
	
	signal bitvectord1906d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1906d : std_logic := '0';
	signal matchd1906d : std_logic := '0';
	
	signal bitvectord1907d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1907d : std_logic := '0';
	signal matchd1907d : std_logic := '0';
	
	signal bitvectord1908d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1908d : std_logic := '0';
	signal matchd1908d : std_logic := '0';
	
	signal bitvectord1909d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1909d : std_logic := '0';
	signal matchd1909d : std_logic := '0';
	
	signal bitvectord1910d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1910d : std_logic := '0';
	signal matchd1910d : std_logic := '0';
	
	signal bitvectord1911d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1911d : std_logic := '0';
	signal matchd1911d : std_logic := '0';
	
	signal bitvectord1912d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1912d : std_logic := '0';
	signal matchd1912d : std_logic := '0';
	
	signal bitvectord1913d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1913d : std_logic := '0';
	signal matchd1913d : std_logic := '0';
	
	signal bitvectord1914d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1914d : std_logic := '0';
	signal matchd1914d : std_logic := '0';
	
	signal bitvectord1915d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1915d : std_logic := '0';
	signal matchd1915d : std_logic := '0';
	
	signal bitvectord1916d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1916d : std_logic := '0';
	signal matchd1916d : std_logic := '0';
	
	signal bitvectord1917d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1917d : std_logic := '1';
	signal matchd1917d : std_logic := '0';
	
	signal bitvectord1918d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1918d : std_logic := '0';
	signal matchd1918d : std_logic := '0';
	
	signal bitvectord1919d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1919d : std_logic := '0';
	signal matchd1919d : std_logic := '0';
	
	signal bitvectord1920d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1920d : std_logic := '0';
	signal matchd1920d : std_logic := '0';
	
	signal bitvectord1921d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1921d : std_logic := '0';
	signal matchd1921d : std_logic := '0';
	
	signal bitvectord1922d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1922d : std_logic := '0';
	signal matchd1922d : std_logic := '0';
	
	signal bitvectord1923d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1923d : std_logic := '0';
	signal matchd1923d : std_logic := '0';
	
	signal bitvectord1924d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1924d : std_logic := '0';
	signal matchd1924d : std_logic := '0';
	
	signal bitvectord1925d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1925d : std_logic := '0';
	signal matchd1925d : std_logic := '0';
	
	signal bitvectord1926d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1926d : std_logic := '0';
	signal matchd1926d : std_logic := '0';
	
	signal bitvectord1927d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1927d : std_logic := '0';
	signal matchd1927d : std_logic := '0';
	
	signal bitvectord1928d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1928d : std_logic := '0';
	signal matchd1928d : std_logic := '0';
	
	signal bitvectord1929d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1929d : std_logic := '0';
	signal matchd1929d : std_logic := '0';
	
	signal bitvectord1930d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1930d : std_logic := '0';
	signal matchd1930d : std_logic := '0';
	
	signal bitvectord1931d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1931d : std_logic := '0';
	signal matchd1931d : std_logic := '0';
	
	signal bitvectord1932d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1932d : std_logic := '0';
	signal matchd1932d : std_logic := '0';
	
	signal bitvectord1933d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1933d : std_logic := '0';
	signal matchd1933d : std_logic := '0';
	
	signal bitvectord1934d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1934d : std_logic := '0';
	signal matchd1934d : std_logic := '0';
	
	signal bitvectord1935d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1935d : std_logic := '1';
	signal matchd1935d : std_logic := '0';
	
	signal bitvectord1936d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1936d : std_logic := '0';
	signal matchd1936d : std_logic := '0';
	
	signal bitvectord1937d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1937d : std_logic := '0';
	signal matchd1937d : std_logic := '0';
	
	signal bitvectord1938d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1938d : std_logic := '0';
	signal matchd1938d : std_logic := '0';
	
	signal bitvectord1939d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1939d : std_logic := '0';
	signal matchd1939d : std_logic := '0';
	
	signal bitvectord1940d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1940d : std_logic := '0';
	signal matchd1940d : std_logic := '0';
	
	signal bitvectord1941d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1941d : std_logic := '0';
	signal matchd1941d : std_logic := '0';
	
	signal bitvectord1942d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1942d : std_logic := '0';
	signal matchd1942d : std_logic := '0';
	
	signal bitvectord1943d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000";
	signal Enabled1943d : std_logic := '0';
	signal matchd1943d : std_logic := '0';
	
	signal bitvectord1944d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1944d : std_logic := '0';
	signal matchd1944d : std_logic := '0';
	
	signal bitvectord1945d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1945d : std_logic := '1';
	signal matchd1945d : std_logic := '0';
	
	signal bitvectord1946d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1946d : std_logic := '0';
	signal matchd1946d : std_logic := '0';
	
	signal bitvectord1947d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1947d : std_logic := '0';
	signal matchd1947d : std_logic := '0';
	
	signal bitvectord1948d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1948d : std_logic := '0';
	signal matchd1948d : std_logic := '0';
	
	signal bitvectord1949d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1949d : std_logic := '0';
	signal matchd1949d : std_logic := '0';
	
	signal bitvectord1950d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1950d : std_logic := '0';
	signal matchd1950d : std_logic := '0';
	
	signal bitvectord1951d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1951d : std_logic := '0';
	signal matchd1951d : std_logic := '0';
	
	signal bitvectord1952d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1952d : std_logic := '0';
	signal matchd1952d : std_logic := '0';
	
	signal bitvectord1953d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1953d : std_logic := '0';
	signal matchd1953d : std_logic := '0';
	
	signal bitvectord1954d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1954d : std_logic := '0';
	signal matchd1954d : std_logic := '0';
	
	signal bitvectord1955d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1955d : std_logic := '0';
	signal matchd1955d : std_logic := '0';
	
	signal bitvectord1956d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1956d : std_logic := '0';
	signal matchd1956d : std_logic := '0';
	
	signal bitvectord1957d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1957d : std_logic := '1';
	signal matchd1957d : std_logic := '0';
	
	signal bitvectord1958d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1958d : std_logic := '0';
	signal matchd1958d : std_logic := '0';
	
	signal bitvectord1959d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1959d : std_logic := '0';
	signal matchd1959d : std_logic := '0';
	
	signal bitvectord1960d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1960d : std_logic := '0';
	signal matchd1960d : std_logic := '0';
	
	signal bitvectord1961d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1961d : std_logic := '0';
	signal matchd1961d : std_logic := '0';
	
	signal bitvectord1962d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1962d : std_logic := '0';
	signal matchd1962d : std_logic := '0';
	
	signal bitvectord1963d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1963d : std_logic := '0';
	signal matchd1963d : std_logic := '0';
	
	signal bitvectord1964d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1964d : std_logic := '0';
	signal matchd1964d : std_logic := '0';
	
	signal bitvectord1965d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1965d : std_logic := '0';
	signal matchd1965d : std_logic := '0';
	
	signal bitvectord1966d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1966d : std_logic := '0';
	signal matchd1966d : std_logic := '0';
	
	signal bitvectord1967d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1967d : std_logic := '0';
	signal matchd1967d : std_logic := '0';
	
	signal bitvectord1968d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1968d : std_logic := '0';
	signal matchd1968d : std_logic := '0';
	
	signal bitvectord1969d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1969d : std_logic := '1';
	signal matchd1969d : std_logic := '0';
	
	signal bitvectord1970d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1970d : std_logic := '0';
	signal matchd1970d : std_logic := '0';
	
	signal bitvectord1971d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1971d : std_logic := '0';
	signal matchd1971d : std_logic := '0';
	
	signal bitvectord1972d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1972d : std_logic := '0';
	signal matchd1972d : std_logic := '0';
	
	signal bitvectord1973d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1973d : std_logic := '0';
	signal matchd1973d : std_logic := '0';
	
	signal bitvectord1974d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1974d : std_logic := '0';
	signal matchd1974d : std_logic := '0';
	
	signal bitvectord1975d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1975d : std_logic := '0';
	signal matchd1975d : std_logic := '0';
	
	signal bitvectord1976d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1976d : std_logic := '0';
	signal matchd1976d : std_logic := '0';
	
	signal bitvectord1977d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1977d : std_logic := '0';
	signal matchd1977d : std_logic := '0';
	
	signal bitvectord1978d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1978d : std_logic := '0';
	signal matchd1978d : std_logic := '0';
	
	signal bitvectord1979d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1979d : std_logic := '0';
	signal matchd1979d : std_logic := '0';
	
	signal bitvectord1980d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1980d : std_logic := '0';
	signal matchd1980d : std_logic := '0';
	
	signal bitvectord1981d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1981d : std_logic := '1';
	signal matchd1981d : std_logic := '0';
	
	signal bitvectord1982d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1982d : std_logic := '0';
	signal matchd1982d : std_logic := '0';
	
	signal bitvectord1983d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1983d : std_logic := '0';
	signal matchd1983d : std_logic := '0';
	
	signal bitvectord1984d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1984d : std_logic := '0';
	signal matchd1984d : std_logic := '0';
	
	signal bitvectord1985d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1985d : std_logic := '0';
	signal matchd1985d : std_logic := '0';
	
	signal bitvectord1986d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1986d : std_logic := '0';
	signal matchd1986d : std_logic := '0';
	
	signal bitvectord1987d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1987d : std_logic := '0';
	signal matchd1987d : std_logic := '0';
	
	signal bitvectord1988d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1988d : std_logic := '0';
	signal matchd1988d : std_logic := '0';
	
	signal bitvectord1989d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1989d : std_logic := '0';
	signal matchd1989d : std_logic := '0';
	
	signal bitvectord1990d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1990d : std_logic := '0';
	signal matchd1990d : std_logic := '0';
	
	signal bitvectord1991d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1991d : std_logic := '0';
	signal matchd1991d : std_logic := '0';
	
	signal bitvectord1992d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1992d : std_logic := '0';
	signal matchd1992d : std_logic := '0';
	
	signal bitvectord1993d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1993d : std_logic := '0';
	signal matchd1993d : std_logic := '0';
	
	signal bitvectord1994d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111";
	signal Enabled1994d : std_logic := '0';
	signal matchd1994d : std_logic := '0';
	
	signal bitvectord1995d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1995d : std_logic := '0';
	signal matchd1995d : std_logic := '0';
	
	signal bitvectord1996d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled1996d : std_logic := '1';
	signal matchd1996d : std_logic := '0';
	
	signal bitvectord1997d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled1997d : std_logic := '0';
	signal matchd1997d : std_logic := '0';
	
	signal bitvectord1998d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled1998d : std_logic := '0';
	signal matchd1998d : std_logic := '0';
	
	signal bitvectord1999d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled1999d : std_logic := '0';
	signal matchd1999d : std_logic := '0';
	
	signal bitvectord2000d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2000d : std_logic := '0';
	signal matchd2000d : std_logic := '0';
	
	signal bitvectord2001d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2001d : std_logic := '0';
	signal matchd2001d : std_logic := '0';
	
	signal bitvectord2002d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2002d : std_logic := '0';
	signal matchd2002d : std_logic := '0';
	
	signal bitvectord2003d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2003d : std_logic := '0';
	signal matchd2003d : std_logic := '0';
	
	signal bitvectord2004d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2004d : std_logic := '0';
	signal matchd2004d : std_logic := '0';
	
	signal bitvectord2005d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2005d : std_logic := '0';
	signal matchd2005d : std_logic := '0';
	
	signal bitvectord2006d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2006d : std_logic := '0';
	signal matchd2006d : std_logic := '0';
	
	signal bitvectord2007d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2007d : std_logic := '0';
	signal matchd2007d : std_logic := '0';
	
	signal bitvectord2008d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2008d : std_logic := '0';
	signal matchd2008d : std_logic := '0';
	
	signal bitvectord2009d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2009d : std_logic := '0';
	signal matchd2009d : std_logic := '0';
	
	signal bitvectord2010d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2010d : std_logic := '0';
	signal matchd2010d : std_logic := '0';
	
	signal bitvectord2011d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2011d : std_logic := '0';
	signal matchd2011d : std_logic := '0';
	
	signal bitvectord2012d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2012d : std_logic := '0';
	signal matchd2012d : std_logic := '0';
	
	signal bitvectord2013d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2013d : std_logic := '0';
	signal matchd2013d : std_logic := '0';
	
	signal bitvectord2014d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2014d : std_logic := '1';
	signal matchd2014d : std_logic := '0';
	
	signal bitvectord2015d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2015d : std_logic := '0';
	signal matchd2015d : std_logic := '0';
	
	signal bitvectord2016d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2016d : std_logic := '0';
	signal matchd2016d : std_logic := '0';
	
	signal bitvectord2017d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2017d : std_logic := '0';
	signal matchd2017d : std_logic := '0';
	
	signal bitvectord2018d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2018d : std_logic := '0';
	signal matchd2018d : std_logic := '0';
	
	signal bitvectord2019d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2019d : std_logic := '0';
	signal matchd2019d : std_logic := '0';
	
	signal bitvectord2020d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2020d : std_logic := '0';
	signal matchd2020d : std_logic := '0';
	
	signal bitvectord2021d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2021d : std_logic := '0';
	signal matchd2021d : std_logic := '0';
	
	signal bitvectord2022d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2022d : std_logic := '0';
	signal matchd2022d : std_logic := '0';
	
	signal bitvectord2023d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2023d : std_logic := '0';
	signal matchd2023d : std_logic := '0';
	
	signal bitvectord2024d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2024d : std_logic := '0';
	signal matchd2024d : std_logic := '0';
	
	signal bitvectord2025d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2025d : std_logic := '0';
	signal matchd2025d : std_logic := '0';
	
	signal bitvectord2026d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2026d : std_logic := '1';
	signal matchd2026d : std_logic := '0';
	
	signal bitvectord2027d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2027d : std_logic := '0';
	signal matchd2027d : std_logic := '0';
	
	signal bitvectord2028d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2028d : std_logic := '0';
	signal matchd2028d : std_logic := '0';
	
	signal bitvectord2029d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2029d : std_logic := '0';
	signal matchd2029d : std_logic := '0';
	
	signal bitvectord2030d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2030d : std_logic := '0';
	signal matchd2030d : std_logic := '0';
	
	signal bitvectord2031d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2031d : std_logic := '0';
	signal matchd2031d : std_logic := '0';
	
	signal bitvectord2032d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2032d : std_logic := '0';
	signal matchd2032d : std_logic := '0';
	
	signal bitvectord2033d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2033d : std_logic := '0';
	signal matchd2033d : std_logic := '0';
	
	signal bitvectord2034d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2034d : std_logic := '0';
	signal matchd2034d : std_logic := '0';
	
	signal bitvectord2035d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2035d : std_logic := '0';
	signal matchd2035d : std_logic := '0';
	
	signal bitvectord2036d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2036d : std_logic := '0';
	signal matchd2036d : std_logic := '0';
	
	signal bitvectord2037d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2037d : std_logic := '0';
	signal matchd2037d : std_logic := '0';
	
	signal bitvectord2038d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2038d : std_logic := '1';
	signal matchd2038d : std_logic := '0';
	
	signal bitvectord2039d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2039d : std_logic := '0';
	signal matchd2039d : std_logic := '0';
	
	signal bitvectord2040d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2040d : std_logic := '0';
	signal matchd2040d : std_logic := '0';
	
	signal bitvectord2041d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2041d : std_logic := '0';
	signal matchd2041d : std_logic := '0';
	
	signal bitvectord2042d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2042d : std_logic := '0';
	signal matchd2042d : std_logic := '0';
	
	signal bitvectord2043d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2043d : std_logic := '0';
	signal matchd2043d : std_logic := '0';
	
	signal bitvectord2044d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2044d : std_logic := '0';
	signal matchd2044d : std_logic := '0';
	
	signal bitvectord2045d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2045d : std_logic := '0';
	signal matchd2045d : std_logic := '0';
	
	signal bitvectord2046d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2046d : std_logic := '0';
	signal matchd2046d : std_logic := '0';
	
	signal bitvectord2047d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2047d : std_logic := '0';
	signal matchd2047d : std_logic := '0';
	
	signal bitvectord2048d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2048d : std_logic := '0';
	signal matchd2048d : std_logic := '0';
	
	signal bitvectord2049d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2049d : std_logic := '0';
	signal matchd2049d : std_logic := '0';
	
	signal bitvectord2050d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2050d : std_logic := '1';
	signal matchd2050d : std_logic := '0';
	
	signal bitvectord2051d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2051d : std_logic := '0';
	signal matchd2051d : std_logic := '0';
	
	signal bitvectord2052d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2052d : std_logic := '0';
	signal matchd2052d : std_logic := '0';
	
	signal bitvectord2053d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2053d : std_logic := '0';
	signal matchd2053d : std_logic := '0';
	
	signal bitvectord2054d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2054d : std_logic := '0';
	signal matchd2054d : std_logic := '0';
	
	signal bitvectord2055d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2055d : std_logic := '0';
	signal matchd2055d : std_logic := '0';
	
	signal bitvectord2056d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2056d : std_logic := '0';
	signal matchd2056d : std_logic := '0';
	
	signal bitvectord2057d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2057d : std_logic := '0';
	signal matchd2057d : std_logic := '0';
	
	signal bitvectord2058d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000";
	signal Enabled2058d : std_logic := '0';
	signal matchd2058d : std_logic := '0';
	
	signal bitvectord2059d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2059d : std_logic := '0';
	signal matchd2059d : std_logic := '0';
	
	signal bitvectord2060d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2060d : std_logic := '0';
	signal matchd2060d : std_logic := '0';
	
	signal bitvectord2061d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2061d : std_logic := '0';
	signal matchd2061d : std_logic := '0';
	
	signal bitvectord2062d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2062d : std_logic := '0';
	signal matchd2062d : std_logic := '0';
	
	signal bitvectord2063d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2063d : std_logic := '0';
	signal matchd2063d : std_logic := '0';
	
	signal bitvectord2064d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2064d : std_logic := '0';
	signal matchd2064d : std_logic := '0';
	
	signal bitvectord2065d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2065d : std_logic := '1';
	signal matchd2065d : std_logic := '0';
	
	signal bitvectord2066d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2066d : std_logic := '0';
	signal matchd2066d : std_logic := '0';
	
	signal bitvectord2067d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2067d : std_logic := '0';
	signal matchd2067d : std_logic := '0';
	
	signal bitvectord2068d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2068d : std_logic := '0';
	signal matchd2068d : std_logic := '0';
	
	signal bitvectord2069d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2069d : std_logic := '0';
	signal matchd2069d : std_logic := '0';
	
	signal bitvectord2070d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2070d : std_logic := '0';
	signal matchd2070d : std_logic := '0';
	
	signal bitvectord2071d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2071d : std_logic := '0';
	signal matchd2071d : std_logic := '0';
	
	signal bitvectord2072d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2072d : std_logic := '0';
	signal matchd2072d : std_logic := '0';
	
	signal bitvectord2073d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2073d : std_logic := '0';
	signal matchd2073d : std_logic := '0';
	
	signal bitvectord2074d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2074d : std_logic := '0';
	signal matchd2074d : std_logic := '0';
	
	signal bitvectord2075d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2075d : std_logic := '0';
	signal matchd2075d : std_logic := '0';
	
	signal bitvectord2076d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2076d : std_logic := '0';
	signal matchd2076d : std_logic := '0';
	
	signal bitvectord2077d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2077d : std_logic := '0';
	signal matchd2077d : std_logic := '0';
	
	signal bitvectord2078d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2078d : std_logic := '0';
	signal matchd2078d : std_logic := '0';
	
	signal bitvectord2079d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2079d : std_logic := '0';
	signal matchd2079d : std_logic := '0';
	
	signal bitvectord2080d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2080d : std_logic := '1';
	signal matchd2080d : std_logic := '0';
	
	signal bitvectord2081d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2081d : std_logic := '0';
	signal matchd2081d : std_logic := '0';
	
	signal bitvectord2082d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2082d : std_logic := '0';
	signal matchd2082d : std_logic := '0';
	
	signal bitvectord2083d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2083d : std_logic := '0';
	signal matchd2083d : std_logic := '0';
	
	signal bitvectord2084d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2084d : std_logic := '0';
	signal matchd2084d : std_logic := '0';
	
	signal bitvectord2085d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2085d : std_logic := '0';
	signal matchd2085d : std_logic := '0';
	
	signal bitvectord2086d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2086d : std_logic := '0';
	signal matchd2086d : std_logic := '0';
	
	signal bitvectord2087d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2087d : std_logic := '0';
	signal matchd2087d : std_logic := '0';
	
	signal bitvectord2088d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2088d : std_logic := '0';
	signal matchd2088d : std_logic := '0';
	
	signal bitvectord2089d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2089d : std_logic := '0';
	signal matchd2089d : std_logic := '0';
	
	signal bitvectord2090d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2090d : std_logic := '0';
	signal matchd2090d : std_logic := '0';
	
	signal bitvectord2091d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2091d : std_logic := '0';
	signal matchd2091d : std_logic := '0';
	
	signal bitvectord2092d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2092d : std_logic := '0';
	signal matchd2092d : std_logic := '0';
	
	signal bitvectord2093d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2093d : std_logic := '0';
	signal matchd2093d : std_logic := '0';
	
	signal bitvectord2094d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2094d : std_logic := '0';
	signal matchd2094d : std_logic := '0';
	
	signal bitvectord2095d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2095d : std_logic := '1';
	signal matchd2095d : std_logic := '0';
	
	signal bitvectord2096d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2096d : std_logic := '0';
	signal matchd2096d : std_logic := '0';
	
	signal bitvectord2097d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2097d : std_logic := '0';
	signal matchd2097d : std_logic := '0';
	
	signal bitvectord2098d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2098d : std_logic := '0';
	signal matchd2098d : std_logic := '0';
	
	signal bitvectord2099d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2099d : std_logic := '0';
	signal matchd2099d : std_logic := '0';
	
	signal bitvectord2100d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2100d : std_logic := '0';
	signal matchd2100d : std_logic := '0';
	
	signal bitvectord2101d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2101d : std_logic := '0';
	signal matchd2101d : std_logic := '0';
	
	signal bitvectord2102d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2102d : std_logic := '0';
	signal matchd2102d : std_logic := '0';
	
	signal bitvectord2103d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2103d : std_logic := '0';
	signal matchd2103d : std_logic := '0';
	
	signal bitvectord2104d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2104d : std_logic := '0';
	signal matchd2104d : std_logic := '0';
	
	signal bitvectord2105d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2105d : std_logic := '0';
	signal matchd2105d : std_logic := '0';
	
	signal bitvectord2106d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2106d : std_logic := '0';
	signal matchd2106d : std_logic := '0';
	
	signal bitvectord2107d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2107d : std_logic := '0';
	signal matchd2107d : std_logic := '0';
	
	signal bitvectord2108d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2108d : std_logic := '1';
	signal matchd2108d : std_logic := '0';
	
	signal bitvectord2109d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2109d : std_logic := '0';
	signal matchd2109d : std_logic := '0';
	
	signal bitvectord2110d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2110d : std_logic := '0';
	signal matchd2110d : std_logic := '0';
	
	signal bitvectord2111d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2111d : std_logic := '0';
	signal matchd2111d : std_logic := '0';
	
	signal bitvectord2112d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2112d : std_logic := '0';
	signal matchd2112d : std_logic := '0';
	
	signal bitvectord2113d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2113d : std_logic := '0';
	signal matchd2113d : std_logic := '0';
	
	signal bitvectord2114d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2114d : std_logic := '0';
	signal matchd2114d : std_logic := '0';
	
	signal bitvectord2115d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2115d : std_logic := '0';
	signal matchd2115d : std_logic := '0';
	
	signal bitvectord2116d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2116d : std_logic := '0';
	signal matchd2116d : std_logic := '0';
	
	signal bitvectord2117d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2117d : std_logic := '0';
	signal matchd2117d : std_logic := '0';
	
	signal bitvectord2118d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2118d : std_logic := '0';
	signal matchd2118d : std_logic := '0';
	
	signal bitvectord2119d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2119d : std_logic := '0';
	signal matchd2119d : std_logic := '0';
	
	signal bitvectord2120d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2120d : std_logic := '1';
	signal matchd2120d : std_logic := '0';
	
	signal bitvectord2121d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2121d : std_logic := '0';
	signal matchd2121d : std_logic := '0';
	
	signal bitvectord2122d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2122d : std_logic := '0';
	signal matchd2122d : std_logic := '0';
	
	signal bitvectord2123d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2123d : std_logic := '0';
	signal matchd2123d : std_logic := '0';
	
	signal bitvectord2124d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2124d : std_logic := '0';
	signal matchd2124d : std_logic := '0';
	
	signal bitvectord2125d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2125d : std_logic := '0';
	signal matchd2125d : std_logic := '0';
	
	signal bitvectord2126d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2126d : std_logic := '0';
	signal matchd2126d : std_logic := '0';
	
	signal bitvectord2127d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2127d : std_logic := '0';
	signal matchd2127d : std_logic := '0';
	
	signal bitvectord2128d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2128d : std_logic := '0';
	signal matchd2128d : std_logic := '0';
	
	signal bitvectord2129d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2129d : std_logic := '0';
	signal matchd2129d : std_logic := '0';
	
	signal bitvectord2130d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2130d : std_logic := '0';
	signal matchd2130d : std_logic := '0';
	
	signal bitvectord2131d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2131d : std_logic := '0';
	signal matchd2131d : std_logic := '0';
	
	signal bitvectord2132d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2132d : std_logic := '0';
	signal matchd2132d : std_logic := '0';
	
	signal bitvectord2133d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2133d : std_logic := '0';
	signal matchd2133d : std_logic := '0';
	
	signal bitvectord2134d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2134d : std_logic := '0';
	signal matchd2134d : std_logic := '0';
	
	signal bitvectord2135d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2135d : std_logic := '0';
	signal matchd2135d : std_logic := '0';
	
	signal bitvectord2136d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2136d : std_logic := '0';
	signal matchd2136d : std_logic := '0';
	
	signal bitvectord2137d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2137d : std_logic := '0';
	signal matchd2137d : std_logic := '0';
	
	signal bitvectord2138d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2138d : std_logic := '0';
	signal matchd2138d : std_logic := '0';
	
	signal bitvectord2139d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2139d : std_logic := '0';
	signal matchd2139d : std_logic := '0';
	
	signal bitvectord2140d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2140d : std_logic := '0';
	signal matchd2140d : std_logic := '0';
	
	signal bitvectord2141d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2141d : std_logic := '0';
	signal matchd2141d : std_logic := '0';
	
	signal bitvectord2142d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2142d : std_logic := '1';
	signal matchd2142d : std_logic := '0';
	
	signal bitvectord2143d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2143d : std_logic := '0';
	signal matchd2143d : std_logic := '0';
	
	signal bitvectord2144d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2144d : std_logic := '0';
	signal matchd2144d : std_logic := '0';
	
	signal bitvectord2145d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2145d : std_logic := '0';
	signal matchd2145d : std_logic := '0';
	
	signal bitvectord2146d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2146d : std_logic := '0';
	signal matchd2146d : std_logic := '0';
	
	signal bitvectord2147d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2147d : std_logic := '0';
	signal matchd2147d : std_logic := '0';
	
	signal bitvectord2148d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2148d : std_logic := '0';
	signal matchd2148d : std_logic := '0';
	
	signal bitvectord2149d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2149d : std_logic := '0';
	signal matchd2149d : std_logic := '0';
	
	signal bitvectord2150d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2150d : std_logic := '0';
	signal matchd2150d : std_logic := '0';
	
	signal bitvectord2151d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2151d : std_logic := '0';
	signal matchd2151d : std_logic := '0';
	
	signal bitvectord2152d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2152d : std_logic := '0';
	signal matchd2152d : std_logic := '0';
	
	signal bitvectord2153d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2153d : std_logic := '0';
	signal matchd2153d : std_logic := '0';
	
	signal bitvectord2154d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2154d : std_logic := '0';
	signal matchd2154d : std_logic := '0';
	
	signal bitvectord2155d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2155d : std_logic := '0';
	signal matchd2155d : std_logic := '0';
	
	signal bitvectord2156d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2156d : std_logic := '0';
	signal matchd2156d : std_logic := '0';
	
	signal bitvectord2157d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2157d : std_logic := '0';
	signal matchd2157d : std_logic := '0';
	
	signal bitvectord2158d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2158d : std_logic := '0';
	signal matchd2158d : std_logic := '0';
	
	signal bitvectord2159d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2159d : std_logic := '1';
	signal matchd2159d : std_logic := '0';
	
	signal bitvectord2160d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2160d : std_logic := '0';
	signal matchd2160d : std_logic := '0';
	
	signal bitvectord2161d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2161d : std_logic := '0';
	signal matchd2161d : std_logic := '0';
	
	signal bitvectord2162d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2162d : std_logic := '0';
	signal matchd2162d : std_logic := '0';
	
	signal bitvectord2163d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2163d : std_logic := '0';
	signal matchd2163d : std_logic := '0';
	
	signal bitvectord2164d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2164d : std_logic := '0';
	signal matchd2164d : std_logic := '0';
	
	signal bitvectord2165d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2165d : std_logic := '0';
	signal matchd2165d : std_logic := '0';
	
	signal bitvectord2166d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2166d : std_logic := '0';
	signal matchd2166d : std_logic := '0';
	
	signal bitvectord2167d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2167d : std_logic := '0';
	signal matchd2167d : std_logic := '0';
	
	signal bitvectord2168d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2168d : std_logic := '0';
	signal matchd2168d : std_logic := '0';
	
	signal bitvectord2169d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2169d : std_logic := '0';
	signal matchd2169d : std_logic := '0';
	
	signal bitvectord2170d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2170d : std_logic := '0';
	signal matchd2170d : std_logic := '0';
	
	signal bitvectord2171d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2171d : std_logic := '1';
	signal matchd2171d : std_logic := '0';
	
	signal bitvectord2172d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2172d : std_logic := '0';
	signal matchd2172d : std_logic := '0';
	
	signal bitvectord2173d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2173d : std_logic := '0';
	signal matchd2173d : std_logic := '0';
	
	signal bitvectord2174d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2174d : std_logic := '0';
	signal matchd2174d : std_logic := '0';
	
	signal bitvectord2175d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2175d : std_logic := '0';
	signal matchd2175d : std_logic := '0';
	
	signal bitvectord2176d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2176d : std_logic := '0';
	signal matchd2176d : std_logic := '0';
	
	signal bitvectord2177d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2177d : std_logic := '0';
	signal matchd2177d : std_logic := '0';
	
	signal bitvectord2178d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2178d : std_logic := '0';
	signal matchd2178d : std_logic := '0';
	
	signal bitvectord2179d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2179d : std_logic := '0';
	signal matchd2179d : std_logic := '0';
	
	signal bitvectord2180d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2180d : std_logic := '0';
	signal matchd2180d : std_logic := '0';
	
	signal bitvectord2181d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2181d : std_logic := '0';
	signal matchd2181d : std_logic := '0';
	
	signal bitvectord2182d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2182d : std_logic := '0';
	signal matchd2182d : std_logic := '0';
	
	signal bitvectord2183d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2183d : std_logic := '0';
	signal matchd2183d : std_logic := '0';
	
	signal bitvectord2184d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2184d : std_logic := '0';
	signal matchd2184d : std_logic := '0';
	
	signal bitvectord2185d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2185d : std_logic := '0';
	signal matchd2185d : std_logic := '0';
	
	signal bitvectord2186d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2186d : std_logic := '0';
	signal matchd2186d : std_logic := '0';
	
	signal bitvectord2187d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2187d : std_logic := '0';
	signal matchd2187d : std_logic := '0';
	
	signal bitvectord2188d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2188d : std_logic := '0';
	signal matchd2188d : std_logic := '0';
	
	signal bitvectord2189d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2189d : std_logic := '0';
	signal matchd2189d : std_logic := '0';
	
	signal bitvectord2190d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2190d : std_logic := '0';
	signal matchd2190d : std_logic := '0';
	
	signal bitvectord2191d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2191d : std_logic := '0';
	signal matchd2191d : std_logic := '0';
	
	signal bitvectord2192d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2192d : std_logic := '0';
	signal matchd2192d : std_logic := '0';
	
	signal bitvectord2193d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2193d : std_logic := '1';
	signal matchd2193d : std_logic := '0';
	
	signal bitvectord2194d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2194d : std_logic := '0';
	signal matchd2194d : std_logic := '0';
	
	signal bitvectord2195d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2195d : std_logic := '0';
	signal matchd2195d : std_logic := '0';
	
	signal bitvectord2196d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2196d : std_logic := '0';
	signal matchd2196d : std_logic := '0';
	
	signal bitvectord2197d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2197d : std_logic := '0';
	signal matchd2197d : std_logic := '0';
	
	signal bitvectord2198d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2198d : std_logic := '0';
	signal matchd2198d : std_logic := '0';
	
	signal bitvectord2199d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2199d : std_logic := '0';
	signal matchd2199d : std_logic := '0';
	
	signal bitvectord2200d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2200d : std_logic := '0';
	signal matchd2200d : std_logic := '0';
	
	signal bitvectord2201d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2201d : std_logic := '0';
	signal matchd2201d : std_logic := '0';
	
	signal bitvectord2202d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2202d : std_logic := '0';
	signal matchd2202d : std_logic := '0';
	
	signal bitvectord2203d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2203d : std_logic := '0';
	signal matchd2203d : std_logic := '0';
	
	signal bitvectord2204d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2204d : std_logic := '0';
	signal matchd2204d : std_logic := '0';
	
	signal bitvectord2205d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2205d : std_logic := '0';
	signal matchd2205d : std_logic := '0';
	
	signal bitvectord2206d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2206d : std_logic := '0';
	signal matchd2206d : std_logic := '0';
	
	signal bitvectord2207d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2207d : std_logic := '0';
	signal matchd2207d : std_logic := '0';
	
	signal bitvectord2208d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2208d : std_logic := '0';
	signal matchd2208d : std_logic := '0';
	
	signal bitvectord2209d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2209d : std_logic := '1';
	signal matchd2209d : std_logic := '0';
	
	signal bitvectord2210d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2210d : std_logic := '0';
	signal matchd2210d : std_logic := '0';
	
	signal bitvectord2211d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2211d : std_logic := '0';
	signal matchd2211d : std_logic := '0';
	
	signal bitvectord2212d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2212d : std_logic := '0';
	signal matchd2212d : std_logic := '0';
	
	signal bitvectord2213d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2213d : std_logic := '0';
	signal matchd2213d : std_logic := '0';
	
	signal bitvectord2214d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2214d : std_logic := '0';
	signal matchd2214d : std_logic := '0';
	
	signal bitvectord2215d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2215d : std_logic := '0';
	signal matchd2215d : std_logic := '0';
	
	signal bitvectord2216d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2216d : std_logic := '0';
	signal matchd2216d : std_logic := '0';
	
	signal bitvectord2217d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2217d : std_logic := '0';
	signal matchd2217d : std_logic := '0';
	
	signal bitvectord2218d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2218d : std_logic := '0';
	signal matchd2218d : std_logic := '0';
	
	signal bitvectord2219d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2219d : std_logic := '0';
	signal matchd2219d : std_logic := '0';
	
	signal bitvectord2220d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2220d : std_logic := '0';
	signal matchd2220d : std_logic := '0';
	
	signal bitvectord2221d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2221d : std_logic := '1';
	signal matchd2221d : std_logic := '0';
	
	signal bitvectord2222d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2222d : std_logic := '0';
	signal matchd2222d : std_logic := '0';
	
	signal bitvectord2223d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2223d : std_logic := '0';
	signal matchd2223d : std_logic := '0';
	
	signal bitvectord2224d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2224d : std_logic := '0';
	signal matchd2224d : std_logic := '0';
	
	signal bitvectord2225d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2225d : std_logic := '0';
	signal matchd2225d : std_logic := '0';
	
	signal bitvectord2226d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2226d : std_logic := '0';
	signal matchd2226d : std_logic := '0';
	
	signal bitvectord2227d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2227d : std_logic := '0';
	signal matchd2227d : std_logic := '0';
	
	signal bitvectord2228d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2228d : std_logic := '0';
	signal matchd2228d : std_logic := '0';
	
	signal bitvectord2229d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2229d : std_logic := '0';
	signal matchd2229d : std_logic := '0';
	
	signal bitvectord2230d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2230d : std_logic := '0';
	signal matchd2230d : std_logic := '0';
	
	signal bitvectord2231d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2231d : std_logic := '0';
	signal matchd2231d : std_logic := '0';
	
	signal bitvectord2232d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2232d : std_logic := '0';
	signal matchd2232d : std_logic := '0';
	
	signal bitvectord2233d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2233d : std_logic := '1';
	signal matchd2233d : std_logic := '0';
	
	signal bitvectord2234d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2234d : std_logic := '0';
	signal matchd2234d : std_logic := '0';
	
	signal bitvectord2235d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2235d : std_logic := '0';
	signal matchd2235d : std_logic := '0';
	
	signal bitvectord2236d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2236d : std_logic := '0';
	signal matchd2236d : std_logic := '0';
	
	signal bitvectord2237d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2237d : std_logic := '0';
	signal matchd2237d : std_logic := '0';
	
	signal bitvectord2238d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2238d : std_logic := '0';
	signal matchd2238d : std_logic := '0';
	
	signal bitvectord2239d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2239d : std_logic := '0';
	signal matchd2239d : std_logic := '0';
	
	signal bitvectord2240d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2240d : std_logic := '0';
	signal matchd2240d : std_logic := '0';
	
	signal bitvectord2241d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2241d : std_logic := '0';
	signal matchd2241d : std_logic := '0';
	
	signal bitvectord2242d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2242d : std_logic := '0';
	signal matchd2242d : std_logic := '0';
	
	signal bitvectord2243d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2243d : std_logic := '0';
	signal matchd2243d : std_logic := '0';
	
	signal bitvectord2244d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2244d : std_logic := '0';
	signal matchd2244d : std_logic := '0';
	
	signal bitvectord2245d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2245d : std_logic := '0';
	signal matchd2245d : std_logic := '0';
	
	signal bitvectord2246d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2246d : std_logic := '0';
	signal matchd2246d : std_logic := '0';
	
	signal bitvectord2247d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2247d : std_logic := '0';
	signal matchd2247d : std_logic := '0';
	
	signal bitvectord2248d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2248d : std_logic := '0';
	signal matchd2248d : std_logic := '0';
	
	signal bitvectord2249d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2249d : std_logic := '0';
	signal matchd2249d : std_logic := '0';
	
	signal bitvectord2250d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000";
	signal Enabled2250d : std_logic := '0';
	signal matchd2250d : std_logic := '0';
	
	signal bitvectord2251d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2251d : std_logic := '0';
	signal matchd2251d : std_logic := '0';
	
	signal bitvectord2252d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2252d : std_logic := '1';
	signal matchd2252d : std_logic := '0';
	
	signal bitvectord2253d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2253d : std_logic := '0';
	signal matchd2253d : std_logic := '0';
	
	signal bitvectord2254d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2254d : std_logic := '0';
	signal matchd2254d : std_logic := '0';
	
	signal bitvectord2255d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2255d : std_logic := '0';
	signal matchd2255d : std_logic := '0';
	
	signal bitvectord2256d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2256d : std_logic := '0';
	signal matchd2256d : std_logic := '0';
	
	signal bitvectord2257d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2257d : std_logic := '0';
	signal matchd2257d : std_logic := '0';
	
	signal bitvectord2258d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2258d : std_logic := '0';
	signal matchd2258d : std_logic := '0';
	
	signal bitvectord2259d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2259d : std_logic := '0';
	signal matchd2259d : std_logic := '0';
	
	signal bitvectord2260d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2260d : std_logic := '0';
	signal matchd2260d : std_logic := '0';
	
	signal bitvectord2261d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2261d : std_logic := '0';
	signal matchd2261d : std_logic := '0';
	
	signal bitvectord2262d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2262d : std_logic := '0';
	signal matchd2262d : std_logic := '0';
	
	signal bitvectord2263d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2263d : std_logic := '0';
	signal matchd2263d : std_logic := '0';
	
	signal bitvectord2264d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2264d : std_logic := '1';
	signal matchd2264d : std_logic := '0';
	
	signal bitvectord2265d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2265d : std_logic := '0';
	signal matchd2265d : std_logic := '0';
	
	signal bitvectord2266d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2266d : std_logic := '0';
	signal matchd2266d : std_logic := '0';
	
	signal bitvectord2267d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2267d : std_logic := '0';
	signal matchd2267d : std_logic := '0';
	
	signal bitvectord2268d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2268d : std_logic := '0';
	signal matchd2268d : std_logic := '0';
	
	signal bitvectord2269d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2269d : std_logic := '0';
	signal matchd2269d : std_logic := '0';
	
	signal bitvectord2270d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2270d : std_logic := '0';
	signal matchd2270d : std_logic := '0';
	
	signal bitvectord2271d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2271d : std_logic := '0';
	signal matchd2271d : std_logic := '0';
	
	signal bitvectord2272d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2272d : std_logic := '0';
	signal matchd2272d : std_logic := '0';
	
	signal bitvectord2273d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2273d : std_logic := '0';
	signal matchd2273d : std_logic := '0';
	
	signal bitvectord2274d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2274d : std_logic := '0';
	signal matchd2274d : std_logic := '0';
	
	signal bitvectord2275d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2275d : std_logic := '0';
	signal matchd2275d : std_logic := '0';
	
	signal bitvectord2276d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2276d : std_logic := '0';
	signal matchd2276d : std_logic := '0';
	
	signal bitvectord2277d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2277d : std_logic := '0';
	signal matchd2277d : std_logic := '0';
	
	signal bitvectord2278d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2278d : std_logic := '0';
	signal matchd2278d : std_logic := '0';
	
	signal bitvectord2279d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2279d : std_logic := '0';
	signal matchd2279d : std_logic := '0';
	
	signal bitvectord2280d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2280d : std_logic := '1';
	signal matchd2280d : std_logic := '0';
	
	signal bitvectord2281d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2281d : std_logic := '0';
	signal matchd2281d : std_logic := '0';
	
	signal bitvectord2282d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2282d : std_logic := '0';
	signal matchd2282d : std_logic := '0';
	
	signal bitvectord2283d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2283d : std_logic := '0';
	signal matchd2283d : std_logic := '0';
	
	signal bitvectord2284d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2284d : std_logic := '0';
	signal matchd2284d : std_logic := '0';
	
	signal bitvectord2285d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2285d : std_logic := '0';
	signal matchd2285d : std_logic := '0';
	
	signal bitvectord2286d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2286d : std_logic := '0';
	signal matchd2286d : std_logic := '0';
	
	signal bitvectord2287d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2287d : std_logic := '0';
	signal matchd2287d : std_logic := '0';
	
	signal bitvectord2288d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2288d : std_logic := '0';
	signal matchd2288d : std_logic := '0';
	
	signal bitvectord2289d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2289d : std_logic := '0';
	signal matchd2289d : std_logic := '0';
	
	signal bitvectord2290d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2290d : std_logic := '0';
	signal matchd2290d : std_logic := '0';
	
	signal bitvectord2291d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2291d : std_logic := '0';
	signal matchd2291d : std_logic := '0';
	
	signal bitvectord2292d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2292d : std_logic := '1';
	signal matchd2292d : std_logic := '0';
	
	signal bitvectord2293d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2293d : std_logic := '0';
	signal matchd2293d : std_logic := '0';
	
	signal bitvectord2294d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2294d : std_logic := '0';
	signal matchd2294d : std_logic := '0';
	
	signal bitvectord2295d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2295d : std_logic := '0';
	signal matchd2295d : std_logic := '0';
	
	signal bitvectord2296d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2296d : std_logic := '0';
	signal matchd2296d : std_logic := '0';
	
	signal bitvectord2297d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2297d : std_logic := '0';
	signal matchd2297d : std_logic := '0';
	
	signal bitvectord2298d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2298d : std_logic := '0';
	signal matchd2298d : std_logic := '0';
	
	signal bitvectord2299d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2299d : std_logic := '0';
	signal matchd2299d : std_logic := '0';
	
	signal bitvectord2300d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2300d : std_logic := '0';
	signal matchd2300d : std_logic := '0';
	
	signal bitvectord2301d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2301d : std_logic := '0';
	signal matchd2301d : std_logic := '0';
	
	signal bitvectord2302d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2302d : std_logic := '0';
	signal matchd2302d : std_logic := '0';
	
	signal bitvectord2303d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2303d : std_logic := '0';
	signal matchd2303d : std_logic := '0';
	
	signal bitvectord2304d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2304d : std_logic := '0';
	signal matchd2304d : std_logic := '0';
	
	signal bitvectord2305d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2305d : std_logic := '0';
	signal matchd2305d : std_logic := '0';
	
	signal bitvectord2306d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2306d : std_logic := '0';
	signal matchd2306d : std_logic := '0';
	
	signal bitvectord2307d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2307d : std_logic := '0';
	signal matchd2307d : std_logic := '0';
	
	signal bitvectord2308d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2308d : std_logic := '1';
	signal matchd2308d : std_logic := '0';
	
	signal bitvectord2309d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2309d : std_logic := '0';
	signal matchd2309d : std_logic := '0';
	
	signal bitvectord2310d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2310d : std_logic := '0';
	signal matchd2310d : std_logic := '0';
	
	signal bitvectord2311d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2311d : std_logic := '0';
	signal matchd2311d : std_logic := '0';
	
	signal bitvectord2312d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2312d : std_logic := '0';
	signal matchd2312d : std_logic := '0';
	
	signal bitvectord2313d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2313d : std_logic := '0';
	signal matchd2313d : std_logic := '0';
	
	signal bitvectord2314d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2314d : std_logic := '0';
	signal matchd2314d : std_logic := '0';
	
	signal bitvectord2315d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2315d : std_logic := '0';
	signal matchd2315d : std_logic := '0';
	
	signal bitvectord2316d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2316d : std_logic := '0';
	signal matchd2316d : std_logic := '0';
	
	signal bitvectord2317d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2317d : std_logic := '0';
	signal matchd2317d : std_logic := '0';
	
	signal bitvectord2318d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2318d : std_logic := '0';
	signal matchd2318d : std_logic := '0';
	
	signal bitvectord2319d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2319d : std_logic := '0';
	signal matchd2319d : std_logic := '0';
	
	signal bitvectord2320d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2320d : std_logic := '0';
	signal matchd2320d : std_logic := '0';
	
	signal bitvectord2321d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2321d : std_logic := '0';
	signal matchd2321d : std_logic := '0';
	
	signal bitvectord2322d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2322d : std_logic := '0';
	signal matchd2322d : std_logic := '0';
	
	signal bitvectord2323d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2323d : std_logic := '0';
	signal matchd2323d : std_logic := '0';
	
	signal bitvectord2325d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2325d : std_logic := '1';
	signal matchd2325d : std_logic := '0';
	
	signal bitvectord2326d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2326d : std_logic := '0';
	signal matchd2326d : std_logic := '0';
	
	signal bitvectord2327d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2327d : std_logic := '0';
	signal matchd2327d : std_logic := '0';
	
	signal bitvectord2328d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2328d : std_logic := '0';
	signal matchd2328d : std_logic := '0';
	
	signal bitvectord2329d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2329d : std_logic := '0';
	signal matchd2329d : std_logic := '0';
	
	signal bitvectord2330d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2330d : std_logic := '0';
	signal matchd2330d : std_logic := '0';
	
	signal bitvectord2331d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2331d : std_logic := '0';
	signal matchd2331d : std_logic := '0';
	
	signal bitvectord2332d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2332d : std_logic := '0';
	signal matchd2332d : std_logic := '0';
	
	signal bitvectord2333d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2333d : std_logic := '0';
	signal matchd2333d : std_logic := '0';
	
	signal bitvectord2334d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2334d : std_logic := '0';
	signal matchd2334d : std_logic := '0';
	
	signal bitvectord2335d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2335d : std_logic := '0';
	signal matchd2335d : std_logic := '0';
	
	signal bitvectord2336d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2336d : std_logic := '0';
	signal matchd2336d : std_logic := '0';
	
	signal bitvectord2337d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2337d : std_logic := '1';
	signal matchd2337d : std_logic := '0';
	
	signal bitvectord2338d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2338d : std_logic := '0';
	signal matchd2338d : std_logic := '0';
	
	signal bitvectord2339d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2339d : std_logic := '0';
	signal matchd2339d : std_logic := '0';
	
	signal bitvectord2340d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2340d : std_logic := '0';
	signal matchd2340d : std_logic := '0';
	
	signal bitvectord2341d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2341d : std_logic := '0';
	signal matchd2341d : std_logic := '0';
	
	signal bitvectord2342d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2342d : std_logic := '0';
	signal matchd2342d : std_logic := '0';
	
	signal bitvectord2343d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2343d : std_logic := '0';
	signal matchd2343d : std_logic := '0';
	
	signal bitvectord2344d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2344d : std_logic := '0';
	signal matchd2344d : std_logic := '0';
	
	signal bitvectord2345d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2345d : std_logic := '0';
	signal matchd2345d : std_logic := '0';
	
	signal bitvectord2346d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2346d : std_logic := '0';
	signal matchd2346d : std_logic := '0';
	
	signal bitvectord2347d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2347d : std_logic := '0';
	signal matchd2347d : std_logic := '0';
	
	signal bitvectord2348d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2348d : std_logic := '0';
	signal matchd2348d : std_logic := '0';
	
	signal bitvectord2349d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2349d : std_logic := '0';
	signal matchd2349d : std_logic := '0';
	
	signal bitvectord2350d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2350d : std_logic := '0';
	signal matchd2350d : std_logic := '0';
	
	signal bitvectord2351d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2351d : std_logic := '0';
	signal matchd2351d : std_logic := '0';
	
	signal bitvectord2352d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2352d : std_logic := '0';
	signal matchd2352d : std_logic := '0';
	
	signal bitvectord2353d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2353d : std_logic := '0';
	signal matchd2353d : std_logic := '0';
	
	signal bitvectord2354d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2354d : std_logic := '1';
	signal matchd2354d : std_logic := '0';
	
	signal bitvectord2355d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2355d : std_logic := '0';
	signal matchd2355d : std_logic := '0';
	
	signal bitvectord2356d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2356d : std_logic := '0';
	signal matchd2356d : std_logic := '0';
	
	signal bitvectord2357d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2357d : std_logic := '0';
	signal matchd2357d : std_logic := '0';
	
	signal bitvectord2358d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2358d : std_logic := '0';
	signal matchd2358d : std_logic := '0';
	
	signal bitvectord2359d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2359d : std_logic := '0';
	signal matchd2359d : std_logic := '0';
	
	signal bitvectord2360d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2360d : std_logic := '0';
	signal matchd2360d : std_logic := '0';
	
	signal bitvectord2361d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2361d : std_logic := '0';
	signal matchd2361d : std_logic := '0';
	
	signal bitvectord2362d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2362d : std_logic := '0';
	signal matchd2362d : std_logic := '0';
	
	signal bitvectord2363d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2363d : std_logic := '0';
	signal matchd2363d : std_logic := '0';
	
	signal bitvectord2364d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2364d : std_logic := '0';
	signal matchd2364d : std_logic := '0';
	
	signal bitvectord2365d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2365d : std_logic := '0';
	signal matchd2365d : std_logic := '0';
	
	signal bitvectord2366d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2366d : std_logic := '0';
	signal matchd2366d : std_logic := '0';
	
	signal bitvectord2367d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2367d : std_logic := '1';
	signal matchd2367d : std_logic := '0';
	
	signal bitvectord2368d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2368d : std_logic := '0';
	signal matchd2368d : std_logic := '0';
	
	signal bitvectord2369d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2369d : std_logic := '0';
	signal matchd2369d : std_logic := '0';
	
	signal bitvectord2370d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2370d : std_logic := '0';
	signal matchd2370d : std_logic := '0';
	
	signal bitvectord2371d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2371d : std_logic := '0';
	signal matchd2371d : std_logic := '0';
	
	signal bitvectord2372d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2372d : std_logic := '0';
	signal matchd2372d : std_logic := '0';
	
	signal bitvectord2373d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2373d : std_logic := '0';
	signal matchd2373d : std_logic := '0';
	
	signal bitvectord2374d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2374d : std_logic := '0';
	signal matchd2374d : std_logic := '0';
	
	signal bitvectord2375d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2375d : std_logic := '0';
	signal matchd2375d : std_logic := '0';
	
	signal bitvectord2376d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2376d : std_logic := '0';
	signal matchd2376d : std_logic := '0';
	
	signal bitvectord2377d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2377d : std_logic := '0';
	signal matchd2377d : std_logic := '0';
	
	signal bitvectord2378d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2378d : std_logic := '0';
	signal matchd2378d : std_logic := '0';
	
	signal bitvectord2379d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2379d : std_logic := '0';
	signal matchd2379d : std_logic := '0';
	
	signal bitvectord2380d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2380d : std_logic := '0';
	signal matchd2380d : std_logic := '0';
	
	signal bitvectord2381d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2381d : std_logic := '0';
	signal matchd2381d : std_logic := '0';
	
	signal bitvectord2382d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2382d : std_logic := '1';
	signal matchd2382d : std_logic := '0';
	
	signal bitvectord2383d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2383d : std_logic := '0';
	signal matchd2383d : std_logic := '0';
	
	signal bitvectord2384d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2384d : std_logic := '0';
	signal matchd2384d : std_logic := '0';
	
	signal bitvectord2385d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2385d : std_logic := '0';
	signal matchd2385d : std_logic := '0';
	
	signal bitvectord2386d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2386d : std_logic := '0';
	signal matchd2386d : std_logic := '0';
	
	signal bitvectord2387d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2387d : std_logic := '0';
	signal matchd2387d : std_logic := '0';
	
	signal bitvectord2388d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2388d : std_logic := '0';
	signal matchd2388d : std_logic := '0';
	
	signal bitvectord2389d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2389d : std_logic := '0';
	signal matchd2389d : std_logic := '0';
	
	signal bitvectord2390d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2390d : std_logic := '0';
	signal matchd2390d : std_logic := '0';
	
	signal bitvectord2391d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2391d : std_logic := '0';
	signal matchd2391d : std_logic := '0';
	
	signal bitvectord2392d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2392d : std_logic := '0';
	signal matchd2392d : std_logic := '0';
	
	signal bitvectord2393d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2393d : std_logic := '0';
	signal matchd2393d : std_logic := '0';
	
	signal bitvectord2394d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2394d : std_logic := '0';
	signal matchd2394d : std_logic := '0';
	
	signal bitvectord2395d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2395d : std_logic := '0';
	signal matchd2395d : std_logic := '0';
	
	signal bitvectord2396d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2396d : std_logic := '0';
	signal matchd2396d : std_logic := '0';
	
	signal bitvectord2398d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2398d : std_logic := '1';
	signal matchd2398d : std_logic := '0';
	
	signal bitvectord2399d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2399d : std_logic := '0';
	signal matchd2399d : std_logic := '0';
	
	signal bitvectord2400d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2400d : std_logic := '0';
	signal matchd2400d : std_logic := '0';
	
	signal bitvectord2401d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2401d : std_logic := '0';
	signal matchd2401d : std_logic := '0';
	
	signal bitvectord2402d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2402d : std_logic := '0';
	signal matchd2402d : std_logic := '0';
	
	signal bitvectord2403d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2403d : std_logic := '0';
	signal matchd2403d : std_logic := '0';
	
	signal bitvectord2404d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2404d : std_logic := '0';
	signal matchd2404d : std_logic := '0';
	
	signal bitvectord2405d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2405d : std_logic := '0';
	signal matchd2405d : std_logic := '0';
	
	signal bitvectord2406d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2406d : std_logic := '0';
	signal matchd2406d : std_logic := '0';
	
	signal bitvectord2407d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2407d : std_logic := '0';
	signal matchd2407d : std_logic := '0';
	
	signal bitvectord2408d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2408d : std_logic := '0';
	signal matchd2408d : std_logic := '0';
	
	signal bitvectord2409d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2409d : std_logic := '0';
	signal matchd2409d : std_logic := '0';
	
	signal bitvectord2410d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2410d : std_logic := '1';
	signal matchd2410d : std_logic := '0';
	
	signal bitvectord2411d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2411d : std_logic := '0';
	signal matchd2411d : std_logic := '0';
	
	signal bitvectord2412d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2412d : std_logic := '0';
	signal matchd2412d : std_logic := '0';
	
	signal bitvectord2413d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2413d : std_logic := '0';
	signal matchd2413d : std_logic := '0';
	
	signal bitvectord2414d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2414d : std_logic := '0';
	signal matchd2414d : std_logic := '0';
	
	signal bitvectord2415d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2415d : std_logic := '0';
	signal matchd2415d : std_logic := '0';
	
	signal bitvectord2416d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2416d : std_logic := '0';
	signal matchd2416d : std_logic := '0';
	
	signal bitvectord2417d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2417d : std_logic := '0';
	signal matchd2417d : std_logic := '0';
	
	signal bitvectord2418d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2418d : std_logic := '0';
	signal matchd2418d : std_logic := '0';
	
	signal bitvectord2419d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2419d : std_logic := '0';
	signal matchd2419d : std_logic := '0';
	
	signal bitvectord2420d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2420d : std_logic := '0';
	signal matchd2420d : std_logic := '0';
	
	signal bitvectord2421d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2421d : std_logic := '1';
	signal matchd2421d : std_logic := '0';
	
	signal bitvectord2422d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2422d : std_logic := '0';
	signal matchd2422d : std_logic := '0';
	
	signal bitvectord2423d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2423d : std_logic := '0';
	signal matchd2423d : std_logic := '0';
	
	signal bitvectord2424d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2424d : std_logic := '0';
	signal matchd2424d : std_logic := '0';
	
	signal bitvectord2425d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2425d : std_logic := '0';
	signal matchd2425d : std_logic := '0';
	
	signal bitvectord2426d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2426d : std_logic := '0';
	signal matchd2426d : std_logic := '0';
	
	signal bitvectord2427d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2427d : std_logic := '0';
	signal matchd2427d : std_logic := '0';
	
	signal bitvectord2428d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2428d : std_logic := '0';
	signal matchd2428d : std_logic := '0';
	
	signal bitvectord2429d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2429d : std_logic := '0';
	signal matchd2429d : std_logic := '0';
	
	signal bitvectord2430d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2430d : std_logic := '0';
	signal matchd2430d : std_logic := '0';
	
	signal bitvectord2431d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2431d : std_logic := '0';
	signal matchd2431d : std_logic := '0';
	
	signal bitvectord2432d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2432d : std_logic := '0';
	signal matchd2432d : std_logic := '0';
	
	signal bitvectord2433d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2433d : std_logic := '0';
	signal matchd2433d : std_logic := '0';
	
	signal bitvectord2434d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2434d : std_logic := '0';
	signal matchd2434d : std_logic := '0';
	
	signal bitvectord2435d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111";
	signal Enabled2435d : std_logic := '0';
	signal matchd2435d : std_logic := '0';
	
	signal bitvectord2436d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2436d : std_logic := '0';
	signal matchd2436d : std_logic := '0';
	
	signal bitvectord2437d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2437d : std_logic := '1';
	signal matchd2437d : std_logic := '0';
	
	signal bitvectord2438d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2438d : std_logic := '0';
	signal matchd2438d : std_logic := '0';
	
	signal bitvectord2439d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2439d : std_logic := '0';
	signal matchd2439d : std_logic := '0';
	
	signal bitvectord2440d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2440d : std_logic := '0';
	signal matchd2440d : std_logic := '0';
	
	signal bitvectord2441d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2441d : std_logic := '0';
	signal matchd2441d : std_logic := '0';
	
	signal bitvectord2442d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2442d : std_logic := '0';
	signal matchd2442d : std_logic := '0';
	
	signal bitvectord2443d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2443d : std_logic := '0';
	signal matchd2443d : std_logic := '0';
	
	signal bitvectord2444d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2444d : std_logic := '0';
	signal matchd2444d : std_logic := '0';
	
	signal bitvectord2445d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2445d : std_logic := '0';
	signal matchd2445d : std_logic := '0';
	
	signal bitvectord2446d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2446d : std_logic := '1';
	signal matchd2446d : std_logic := '0';
	
	signal bitvectord2447d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2447d : std_logic := '0';
	signal matchd2447d : std_logic := '0';
	
	signal bitvectord2448d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2448d : std_logic := '0';
	signal matchd2448d : std_logic := '0';
	
	signal bitvectord2449d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2449d : std_logic := '0';
	signal matchd2449d : std_logic := '0';
	
	signal bitvectord2450d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2450d : std_logic := '0';
	signal matchd2450d : std_logic := '0';
	
	signal bitvectord2451d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2451d : std_logic := '0';
	signal matchd2451d : std_logic := '0';
	
	signal bitvectord2452d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2452d : std_logic := '0';
	signal matchd2452d : std_logic := '0';
	
	signal bitvectord2453d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2453d : std_logic := '0';
	signal matchd2453d : std_logic := '0';
	
	signal bitvectord2454d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2454d : std_logic := '0';
	signal matchd2454d : std_logic := '0';
	
	signal bitvectord2455d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2455d : std_logic := '0';
	signal matchd2455d : std_logic := '0';
	
	signal bitvectord2456d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2456d : std_logic := '0';
	signal matchd2456d : std_logic := '0';
	
	signal bitvectord2457d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2457d : std_logic := '0';
	signal matchd2457d : std_logic := '0';
	
	signal bitvectord2458d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2458d : std_logic := '0';
	signal matchd2458d : std_logic := '0';
	
	signal bitvectord2459d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2459d : std_logic := '0';
	signal matchd2459d : std_logic := '0';
	
	signal bitvectord2460d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2460d : std_logic := '0';
	signal matchd2460d : std_logic := '0';
	
	signal bitvectord2461d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2461d : std_logic := '1';
	signal matchd2461d : std_logic := '0';
	
	signal bitvectord2462d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2462d : std_logic := '0';
	signal matchd2462d : std_logic := '0';
	
	signal bitvectord2463d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2463d : std_logic := '0';
	signal matchd2463d : std_logic := '0';
	
	signal bitvectord2464d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2464d : std_logic := '0';
	signal matchd2464d : std_logic := '0';
	
	signal bitvectord2465d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2465d : std_logic := '0';
	signal matchd2465d : std_logic := '0';
	
	signal bitvectord2466d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2466d : std_logic := '0';
	signal matchd2466d : std_logic := '0';
	
	signal bitvectord2467d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2467d : std_logic := '0';
	signal matchd2467d : std_logic := '0';
	
	signal bitvectord2468d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2468d : std_logic := '0';
	signal matchd2468d : std_logic := '0';
	
	signal bitvectord2469d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2469d : std_logic := '0';
	signal matchd2469d : std_logic := '0';
	
	signal bitvectord2470d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2470d : std_logic := '0';
	signal matchd2470d : std_logic := '0';
	
	signal bitvectord2471d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2471d : std_logic := '0';
	signal matchd2471d : std_logic := '0';
	
	signal bitvectord2472d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2472d : std_logic := '0';
	signal matchd2472d : std_logic := '0';
	
	signal bitvectord2473d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2473d : std_logic := '1';
	signal matchd2473d : std_logic := '0';
	
	signal bitvectord2474d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2474d : std_logic := '0';
	signal matchd2474d : std_logic := '0';
	
	signal bitvectord2475d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2475d : std_logic := '0';
	signal matchd2475d : std_logic := '0';
	
	signal bitvectord2476d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2476d : std_logic := '0';
	signal matchd2476d : std_logic := '0';
	
	signal bitvectord2477d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2477d : std_logic := '0';
	signal matchd2477d : std_logic := '0';
	
	signal bitvectord2478d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2478d : std_logic := '0';
	signal matchd2478d : std_logic := '0';
	
	signal bitvectord2479d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2479d : std_logic := '0';
	signal matchd2479d : std_logic := '0';
	
	signal bitvectord2480d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2480d : std_logic := '0';
	signal matchd2480d : std_logic := '0';
	
	signal bitvectord2481d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2481d : std_logic := '0';
	signal matchd2481d : std_logic := '0';
	
	signal bitvectord2482d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2482d : std_logic := '0';
	signal matchd2482d : std_logic := '0';
	
	signal bitvectord2483d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2483d : std_logic := '0';
	signal matchd2483d : std_logic := '0';
	
	signal bitvectord2484d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2484d : std_logic := '1';
	signal matchd2484d : std_logic := '0';
	
	signal bitvectord2485d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2485d : std_logic := '0';
	signal matchd2485d : std_logic := '0';
	
	signal bitvectord2486d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2486d : std_logic := '0';
	signal matchd2486d : std_logic := '0';
	
	signal bitvectord2487d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2487d : std_logic := '0';
	signal matchd2487d : std_logic := '0';
	
	signal bitvectord2488d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2488d : std_logic := '0';
	signal matchd2488d : std_logic := '0';
	
	signal bitvectord2489d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2489d : std_logic := '0';
	signal matchd2489d : std_logic := '0';
	
	signal bitvectord2490d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2490d : std_logic := '0';
	signal matchd2490d : std_logic := '0';
	
	signal bitvectord2491d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2491d : std_logic := '0';
	signal matchd2491d : std_logic := '0';
	
	signal bitvectord2492d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2492d : std_logic := '0';
	signal matchd2492d : std_logic := '0';
	
	signal bitvectord2493d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2493d : std_logic := '0';
	signal matchd2493d : std_logic := '0';
	
	signal bitvectord2494d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2494d : std_logic := '0';
	signal matchd2494d : std_logic := '0';
	
	signal bitvectord2495d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2495d : std_logic := '0';
	signal matchd2495d : std_logic := '0';
	
	signal bitvectord2496d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2496d : std_logic := '0';
	signal matchd2496d : std_logic := '0';
	
	signal bitvectord2497d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2497d : std_logic := '0';
	signal matchd2497d : std_logic := '0';
	
	signal bitvectord2498d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2498d : std_logic := '0';
	signal matchd2498d : std_logic := '0';
	
	signal bitvectord2499d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2499d : std_logic := '0';
	signal matchd2499d : std_logic := '0';
	
	signal bitvectord2500d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2500d : std_logic := '1';
	signal matchd2500d : std_logic := '0';
	
	signal bitvectord2501d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2501d : std_logic := '0';
	signal matchd2501d : std_logic := '0';
	
	signal bitvectord2502d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2502d : std_logic := '0';
	signal matchd2502d : std_logic := '0';
	
	signal bitvectord2503d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2503d : std_logic := '0';
	signal matchd2503d : std_logic := '0';
	
	signal bitvectord2504d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2504d : std_logic := '0';
	signal matchd2504d : std_logic := '0';
	
	signal bitvectord2505d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2505d : std_logic := '0';
	signal matchd2505d : std_logic := '0';
	
	signal bitvectord2506d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2506d : std_logic := '0';
	signal matchd2506d : std_logic := '0';
	
	signal bitvectord2507d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2507d : std_logic := '0';
	signal matchd2507d : std_logic := '0';
	
	signal bitvectord2508d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2508d : std_logic := '0';
	signal matchd2508d : std_logic := '0';
	
	signal bitvectord2509d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2509d : std_logic := '0';
	signal matchd2509d : std_logic := '0';
	
	signal bitvectord2510d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2510d : std_logic := '0';
	signal matchd2510d : std_logic := '0';
	
	signal bitvectord2511d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2511d : std_logic := '0';
	signal matchd2511d : std_logic := '0';
	
	signal bitvectord2512d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2512d : std_logic := '0';
	signal matchd2512d : std_logic := '0';
	
	signal bitvectord2513d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2513d : std_logic := '0';
	signal matchd2513d : std_logic := '0';
	
	signal bitvectord2514d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2514d : std_logic := '0';
	signal matchd2514d : std_logic := '0';
	
	signal bitvectord2515d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2515d : std_logic := '0';
	signal matchd2515d : std_logic := '0';
	
	signal bitvectord2516d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2516d : std_logic := '0';
	signal matchd2516d : std_logic := '0';
	
	signal bitvectord2517d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2517d : std_logic := '0';
	signal matchd2517d : std_logic := '0';
	
	signal bitvectord2518d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2518d : std_logic := '0';
	signal matchd2518d : std_logic := '0';
	
	signal bitvectord2519d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2519d : std_logic := '0';
	signal matchd2519d : std_logic := '0';
	
	signal bitvectord2520d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2520d : std_logic := '0';
	signal matchd2520d : std_logic := '0';
	
	signal bitvectord2521d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2521d : std_logic := '1';
	signal matchd2521d : std_logic := '0';
	
	signal bitvectord2522d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2522d : std_logic := '0';
	signal matchd2522d : std_logic := '0';
	
	signal bitvectord2523d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2523d : std_logic := '0';
	signal matchd2523d : std_logic := '0';
	
	signal bitvectord2524d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2524d : std_logic := '0';
	signal matchd2524d : std_logic := '0';
	
	signal bitvectord2525d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2525d : std_logic := '0';
	signal matchd2525d : std_logic := '0';
	
	signal bitvectord2526d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2526d : std_logic := '0';
	signal matchd2526d : std_logic := '0';
	
	signal bitvectord2527d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2527d : std_logic := '0';
	signal matchd2527d : std_logic := '0';
	
	signal bitvectord2528d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2528d : std_logic := '0';
	signal matchd2528d : std_logic := '0';
	
	signal bitvectord2529d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2529d : std_logic := '0';
	signal matchd2529d : std_logic := '0';
	
	signal bitvectord2530d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2530d : std_logic := '0';
	signal matchd2530d : std_logic := '0';
	
	signal bitvectord2531d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2531d : std_logic := '0';
	signal matchd2531d : std_logic := '0';
	
	signal bitvectord2532d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2532d : std_logic := '0';
	signal matchd2532d : std_logic := '0';
	
	signal bitvectord2533d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2533d : std_logic := '1';
	signal matchd2533d : std_logic := '0';
	
	signal bitvectord2534d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2534d : std_logic := '0';
	signal matchd2534d : std_logic := '0';
	
	signal bitvectord2535d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2535d : std_logic := '0';
	signal matchd2535d : std_logic := '0';
	
	signal bitvectord2536d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2536d : std_logic := '0';
	signal matchd2536d : std_logic := '0';
	
	signal bitvectord2537d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2537d : std_logic := '0';
	signal matchd2537d : std_logic := '0';
	
	signal bitvectord2538d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2538d : std_logic := '0';
	signal matchd2538d : std_logic := '0';
	
	signal bitvectord2539d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2539d : std_logic := '0';
	signal matchd2539d : std_logic := '0';
	
	signal bitvectord2540d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2540d : std_logic := '0';
	signal matchd2540d : std_logic := '0';
	
	signal bitvectord2541d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2541d : std_logic := '0';
	signal matchd2541d : std_logic := '0';
	
	signal bitvectord2542d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2542d : std_logic := '0';
	signal matchd2542d : std_logic := '0';
	
	signal bitvectord2543d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2543d : std_logic := '0';
	signal matchd2543d : std_logic := '0';
	
	signal bitvectord2544d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2544d : std_logic := '0';
	signal matchd2544d : std_logic := '0';
	
	signal bitvectord2545d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2545d : std_logic := '1';
	signal matchd2545d : std_logic := '0';
	
	signal bitvectord2546d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2546d : std_logic := '0';
	signal matchd2546d : std_logic := '0';
	
	signal bitvectord2547d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2547d : std_logic := '0';
	signal matchd2547d : std_logic := '0';
	
	signal bitvectord2548d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2548d : std_logic := '0';
	signal matchd2548d : std_logic := '0';
	
	signal bitvectord2549d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2549d : std_logic := '0';
	signal matchd2549d : std_logic := '0';
	
	signal bitvectord2550d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2550d : std_logic := '0';
	signal matchd2550d : std_logic := '0';
	
	signal bitvectord2551d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2551d : std_logic := '0';
	signal matchd2551d : std_logic := '0';
	
	signal bitvectord2552d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2552d : std_logic := '0';
	signal matchd2552d : std_logic := '0';
	
	signal bitvectord2553d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2553d : std_logic := '0';
	signal matchd2553d : std_logic := '0';
	
	signal bitvectord2554d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2554d : std_logic := '0';
	signal matchd2554d : std_logic := '0';
	
	signal bitvectord2555d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2555d : std_logic := '0';
	signal matchd2555d : std_logic := '0';
	
	signal bitvectord2556d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2556d : std_logic := '0';
	signal matchd2556d : std_logic := '0';
	
	signal bitvectord2557d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2557d : std_logic := '0';
	signal matchd2557d : std_logic := '0';
	
	signal bitvectord2558d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2558d : std_logic := '0';
	signal matchd2558d : std_logic := '0';
	
	signal bitvectord2559d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2559d : std_logic := '0';
	signal matchd2559d : std_logic := '0';
	
	signal bitvectord2560d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2560d : std_logic := '0';
	signal matchd2560d : std_logic := '0';
	
	signal bitvectord2561d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2561d : std_logic := '0';
	signal matchd2561d : std_logic := '0';
	
	signal bitvectord2562d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2562d : std_logic := '1';
	signal matchd2562d : std_logic := '0';
	
	signal bitvectord2563d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2563d : std_logic := '0';
	signal matchd2563d : std_logic := '0';
	
	signal bitvectord2564d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2564d : std_logic := '0';
	signal matchd2564d : std_logic := '0';
	
	signal bitvectord2565d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2565d : std_logic := '0';
	signal matchd2565d : std_logic := '0';
	
	signal bitvectord2566d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2566d : std_logic := '0';
	signal matchd2566d : std_logic := '0';
	
	signal bitvectord2567d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2567d : std_logic := '0';
	signal matchd2567d : std_logic := '0';
	
	signal bitvectord2568d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2568d : std_logic := '0';
	signal matchd2568d : std_logic := '0';
	
	signal bitvectord2569d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2569d : std_logic := '0';
	signal matchd2569d : std_logic := '0';
	
	signal bitvectord2570d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2570d : std_logic := '0';
	signal matchd2570d : std_logic := '0';
	
	signal bitvectord2571d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2571d : std_logic := '0';
	signal matchd2571d : std_logic := '0';
	
	signal bitvectord2572d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2572d : std_logic := '0';
	signal matchd2572d : std_logic := '0';
	
	signal bitvectord2573d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2573d : std_logic := '1';
	signal matchd2573d : std_logic := '0';
	
	signal bitvectord2574d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2574d : std_logic := '0';
	signal matchd2574d : std_logic := '0';
	
	signal bitvectord2575d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2575d : std_logic := '0';
	signal matchd2575d : std_logic := '0';
	
	signal bitvectord2576d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2576d : std_logic := '0';
	signal matchd2576d : std_logic := '0';
	
	signal bitvectord2577d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2577d : std_logic := '0';
	signal matchd2577d : std_logic := '0';
	
	signal bitvectord2578d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2578d : std_logic := '0';
	signal matchd2578d : std_logic := '0';
	
	signal bitvectord2579d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2579d : std_logic := '0';
	signal matchd2579d : std_logic := '0';
	
	signal bitvectord2580d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2580d : std_logic := '0';
	signal matchd2580d : std_logic := '0';
	
	signal bitvectord2581d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2581d : std_logic := '0';
	signal matchd2581d : std_logic := '0';
	
	signal bitvectord2582d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2582d : std_logic := '0';
	signal matchd2582d : std_logic := '0';
	
	signal bitvectord2583d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2583d : std_logic := '0';
	signal matchd2583d : std_logic := '0';
	
	signal bitvectord2584d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2584d : std_logic := '0';
	signal matchd2584d : std_logic := '0';
	
	signal bitvectord2585d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2585d : std_logic := '0';
	signal matchd2585d : std_logic := '0';
	
	signal bitvectord2586d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2586d : std_logic := '0';
	signal matchd2586d : std_logic := '0';
	
	signal bitvectord2587d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2587d : std_logic := '0';
	signal matchd2587d : std_logic := '0';
	
	signal bitvectord2588d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2588d : std_logic := '0';
	signal matchd2588d : std_logic := '0';
	
	signal bitvectord2589d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2589d : std_logic := '1';
	signal matchd2589d : std_logic := '0';
	
	signal bitvectord2590d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2590d : std_logic := '0';
	signal matchd2590d : std_logic := '0';
	
	signal bitvectord2591d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2591d : std_logic := '0';
	signal matchd2591d : std_logic := '0';
	
	signal bitvectord2592d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2592d : std_logic := '0';
	signal matchd2592d : std_logic := '0';
	
	signal bitvectord2593d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2593d : std_logic := '0';
	signal matchd2593d : std_logic := '0';
	
	signal bitvectord2594d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2594d : std_logic := '0';
	signal matchd2594d : std_logic := '0';
	
	signal bitvectord2595d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2595d : std_logic := '0';
	signal matchd2595d : std_logic := '0';
	
	signal bitvectord2596d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2596d : std_logic := '0';
	signal matchd2596d : std_logic := '0';
	
	signal bitvectord2597d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2597d : std_logic := '0';
	signal matchd2597d : std_logic := '0';
	
	signal bitvectord2598d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2598d : std_logic := '0';
	signal matchd2598d : std_logic := '0';
	
	signal bitvectord2599d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2599d : std_logic := '0';
	signal matchd2599d : std_logic := '0';
	
	signal bitvectord2600d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2600d : std_logic := '1';
	signal matchd2600d : std_logic := '0';
	
	signal bitvectord2601d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2601d : std_logic := '0';
	signal matchd2601d : std_logic := '0';
	
	signal bitvectord2602d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2602d : std_logic := '0';
	signal matchd2602d : std_logic := '0';
	
	signal bitvectord2603d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2603d : std_logic := '0';
	signal matchd2603d : std_logic := '0';
	
	signal bitvectord2604d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2604d : std_logic := '0';
	signal matchd2604d : std_logic := '0';
	
	signal bitvectord2605d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2605d : std_logic := '0';
	signal matchd2605d : std_logic := '0';
	
	signal bitvectord2606d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2606d : std_logic := '0';
	signal matchd2606d : std_logic := '0';
	
	signal bitvectord2607d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2607d : std_logic := '0';
	signal matchd2607d : std_logic := '0';
	
	signal bitvectord2608d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2608d : std_logic := '0';
	signal matchd2608d : std_logic := '0';
	
	signal bitvectord2609d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2609d : std_logic := '0';
	signal matchd2609d : std_logic := '0';
	
	signal bitvectord2610d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2610d : std_logic := '0';
	signal matchd2610d : std_logic := '0';
	
	signal bitvectord2611d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2611d : std_logic := '0';
	signal matchd2611d : std_logic := '0';
	
	signal bitvectord2612d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2612d : std_logic := '0';
	signal matchd2612d : std_logic := '0';
	
	signal bitvectord2613d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2613d : std_logic := '0';
	signal matchd2613d : std_logic := '0';
	
	signal bitvectord2614d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2614d : std_logic := '0';
	signal matchd2614d : std_logic := '0';
	
	signal bitvectord2615d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2615d : std_logic := '0';
	signal matchd2615d : std_logic := '0';
	
	signal bitvectord2616d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2616d : std_logic := '0';
	signal matchd2616d : std_logic := '0';
	
	signal bitvectord2617d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2617d : std_logic := '0';
	signal matchd2617d : std_logic := '0';
	
	signal bitvectord2618d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2618d : std_logic := '0';
	signal matchd2618d : std_logic := '0';
	
	signal bitvectord2619d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2619d : std_logic := '1';
	signal matchd2619d : std_logic := '0';
	
	signal bitvectord2620d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2620d : std_logic := '0';
	signal matchd2620d : std_logic := '0';
	
	signal bitvectord2621d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2621d : std_logic := '0';
	signal matchd2621d : std_logic := '0';
	
	signal bitvectord2622d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2622d : std_logic := '0';
	signal matchd2622d : std_logic := '0';
	
	signal bitvectord2623d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2623d : std_logic := '0';
	signal matchd2623d : std_logic := '0';
	
	signal bitvectord2624d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2624d : std_logic := '0';
	signal matchd2624d : std_logic := '0';
	
	signal bitvectord2625d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2625d : std_logic := '0';
	signal matchd2625d : std_logic := '0';
	
	signal bitvectord2626d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2626d : std_logic := '0';
	signal matchd2626d : std_logic := '0';
	
	signal bitvectord2627d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2627d : std_logic := '0';
	signal matchd2627d : std_logic := '0';
	
	signal bitvectord2628d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2628d : std_logic := '0';
	signal matchd2628d : std_logic := '0';
	
	signal bitvectord2629d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2629d : std_logic := '0';
	signal matchd2629d : std_logic := '0';
	
	signal bitvectord2630d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2630d : std_logic := '0';
	signal matchd2630d : std_logic := '0';
	
	signal bitvectord2631d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2631d : std_logic := '0';
	signal matchd2631d : std_logic := '0';
	
	signal bitvectord2632d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2632d : std_logic := '0';
	signal matchd2632d : std_logic := '0';
	
	signal bitvectord2633d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2633d : std_logic := '0';
	signal matchd2633d : std_logic := '0';
	
	signal bitvectord2634d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000";
	signal Enabled2634d : std_logic := '0';
	signal matchd2634d : std_logic := '0';
	
	signal bitvectord2635d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2635d : std_logic := '0';
	signal matchd2635d : std_logic := '0';
	
	signal bitvectord2636d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2636d : std_logic := '1';
	signal matchd2636d : std_logic := '0';
	
	signal bitvectord2637d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2637d : std_logic := '0';
	signal matchd2637d : std_logic := '0';
	
	signal bitvectord2638d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2638d : std_logic := '0';
	signal matchd2638d : std_logic := '0';
	
	signal bitvectord2639d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2639d : std_logic := '0';
	signal matchd2639d : std_logic := '0';
	
	signal bitvectord2640d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2640d : std_logic := '0';
	signal matchd2640d : std_logic := '0';
	
	signal bitvectord2641d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2641d : std_logic := '0';
	signal matchd2641d : std_logic := '0';
	
	signal bitvectord2642d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2642d : std_logic := '0';
	signal matchd2642d : std_logic := '0';
	
	signal bitvectord2643d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2643d : std_logic := '0';
	signal matchd2643d : std_logic := '0';
	
	signal bitvectord2644d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2644d : std_logic := '0';
	signal matchd2644d : std_logic := '0';
	
	signal bitvectord2645d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2645d : std_logic := '0';
	signal matchd2645d : std_logic := '0';
	
	signal bitvectord2646d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2646d : std_logic := '0';
	signal matchd2646d : std_logic := '0';
	
	signal bitvectord2647d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2647d : std_logic := '0';
	signal matchd2647d : std_logic := '0';
	
	signal bitvectord2648d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2648d : std_logic := '1';
	signal matchd2648d : std_logic := '0';
	
	signal bitvectord2649d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2649d : std_logic := '0';
	signal matchd2649d : std_logic := '0';
	
	signal bitvectord2650d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2650d : std_logic := '0';
	signal matchd2650d : std_logic := '0';
	
	signal bitvectord2651d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2651d : std_logic := '0';
	signal matchd2651d : std_logic := '0';
	
	signal bitvectord2652d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2652d : std_logic := '0';
	signal matchd2652d : std_logic := '0';
	
	signal bitvectord2653d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2653d : std_logic := '0';
	signal matchd2653d : std_logic := '0';
	
	signal bitvectord2654d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2654d : std_logic := '0';
	signal matchd2654d : std_logic := '0';
	
	signal bitvectord2655d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2655d : std_logic := '0';
	signal matchd2655d : std_logic := '0';
	
	signal bitvectord2656d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2656d : std_logic := '0';
	signal matchd2656d : std_logic := '0';
	
	signal bitvectord2657d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2657d : std_logic := '0';
	signal matchd2657d : std_logic := '0';
	
	signal bitvectord2658d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2658d : std_logic := '0';
	signal matchd2658d : std_logic := '0';
	
	signal bitvectord2659d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2659d : std_logic := '0';
	signal matchd2659d : std_logic := '0';
	
	signal bitvectord2660d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2660d : std_logic := '1';
	signal matchd2660d : std_logic := '0';
	
	signal bitvectord2661d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2661d : std_logic := '0';
	signal matchd2661d : std_logic := '0';
	
	signal bitvectord2662d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2662d : std_logic := '0';
	signal matchd2662d : std_logic := '0';
	
	signal bitvectord2663d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2663d : std_logic := '0';
	signal matchd2663d : std_logic := '0';
	
	signal bitvectord2664d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2664d : std_logic := '0';
	signal matchd2664d : std_logic := '0';
	
	signal bitvectord2665d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2665d : std_logic := '0';
	signal matchd2665d : std_logic := '0';
	
	signal bitvectord2666d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2666d : std_logic := '0';
	signal matchd2666d : std_logic := '0';
	
	signal bitvectord2667d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2667d : std_logic := '0';
	signal matchd2667d : std_logic := '0';
	
	signal bitvectord2668d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2668d : std_logic := '0';
	signal matchd2668d : std_logic := '0';
	
	signal bitvectord2669d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2669d : std_logic := '0';
	signal matchd2669d : std_logic := '0';
	
	signal bitvectord2670d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2670d : std_logic := '0';
	signal matchd2670d : std_logic := '0';
	
	signal bitvectord2671d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2671d : std_logic := '0';
	signal matchd2671d : std_logic := '0';
	
	signal bitvectord2672d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2672d : std_logic := '1';
	signal matchd2672d : std_logic := '0';
	
	signal bitvectord2673d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2673d : std_logic := '0';
	signal matchd2673d : std_logic := '0';
	
	signal bitvectord2674d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2674d : std_logic := '0';
	signal matchd2674d : std_logic := '0';
	
	signal bitvectord2675d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2675d : std_logic := '0';
	signal matchd2675d : std_logic := '0';
	
	signal bitvectord2676d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2676d : std_logic := '0';
	signal matchd2676d : std_logic := '0';
	
	signal bitvectord2677d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2677d : std_logic := '0';
	signal matchd2677d : std_logic := '0';
	
	signal bitvectord2678d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2678d : std_logic := '0';
	signal matchd2678d : std_logic := '0';
	
	signal bitvectord2679d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2679d : std_logic := '0';
	signal matchd2679d : std_logic := '0';
	
	signal bitvectord2680d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2680d : std_logic := '0';
	signal matchd2680d : std_logic := '0';
	
	signal bitvectord2681d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2681d : std_logic := '0';
	signal matchd2681d : std_logic := '0';
	
	signal bitvectord2682d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2682d : std_logic := '0';
	signal matchd2682d : std_logic := '0';
	
	signal bitvectord2683d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2683d : std_logic := '0';
	signal matchd2683d : std_logic := '0';
	
	signal bitvectord2684d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2684d : std_logic := '0';
	signal matchd2684d : std_logic := '0';
	
	signal bitvectord2685d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2685d : std_logic := '0';
	signal matchd2685d : std_logic := '0';
	
	signal bitvectord2686d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2686d : std_logic := '0';
	signal matchd2686d : std_logic := '0';
	
	signal bitvectord2687d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2687d : std_logic := '0';
	signal matchd2687d : std_logic := '0';
	
	signal bitvectord2688d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2688d : std_logic := '1';
	signal matchd2688d : std_logic := '0';
	
	signal bitvectord2689d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2689d : std_logic := '0';
	signal matchd2689d : std_logic := '0';
	
	signal bitvectord2690d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2690d : std_logic := '0';
	signal matchd2690d : std_logic := '0';
	
	signal bitvectord2691d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2691d : std_logic := '0';
	signal matchd2691d : std_logic := '0';
	
	signal bitvectord2692d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2692d : std_logic := '0';
	signal matchd2692d : std_logic := '0';
	
	signal bitvectord2693d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2693d : std_logic := '0';
	signal matchd2693d : std_logic := '0';
	
	signal bitvectord2694d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2694d : std_logic := '0';
	signal matchd2694d : std_logic := '0';
	
	signal bitvectord2695d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2695d : std_logic := '0';
	signal matchd2695d : std_logic := '0';
	
	signal bitvectord2696d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2696d : std_logic := '0';
	signal matchd2696d : std_logic := '0';
	
	signal bitvectord2697d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2697d : std_logic := '0';
	signal matchd2697d : std_logic := '0';
	
	signal bitvectord2698d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2698d : std_logic := '1';
	signal matchd2698d : std_logic := '0';
	
	signal bitvectord2699d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2699d : std_logic := '0';
	signal matchd2699d : std_logic := '0';
	
	signal bitvectord2700d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2700d : std_logic := '0';
	signal matchd2700d : std_logic := '0';
	
	signal bitvectord2701d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2701d : std_logic := '0';
	signal matchd2701d : std_logic := '0';
	
	signal bitvectord2702d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2702d : std_logic := '0';
	signal matchd2702d : std_logic := '0';
	
	signal bitvectord2703d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2703d : std_logic := '0';
	signal matchd2703d : std_logic := '0';
	
	signal bitvectord2704d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2704d : std_logic := '0';
	signal matchd2704d : std_logic := '0';
	
	signal bitvectord2705d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2705d : std_logic := '0';
	signal matchd2705d : std_logic := '0';
	
	signal bitvectord2706d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2706d : std_logic := '0';
	signal matchd2706d : std_logic := '0';
	
	signal bitvectord2707d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2707d : std_logic := '0';
	signal matchd2707d : std_logic := '0';
	
	signal bitvectord2708d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2708d : std_logic := '0';
	signal matchd2708d : std_logic := '0';
	
	signal bitvectord2709d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2709d : std_logic := '0';
	signal matchd2709d : std_logic := '0';
	
	signal bitvectord2710d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2710d : std_logic := '0';
	signal matchd2710d : std_logic := '0';
	
	signal bitvectord2711d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000";
	signal Enabled2711d : std_logic := '0';
	signal matchd2711d : std_logic := '0';
	
	signal bitvectord2712d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2712d : std_logic := '0';
	signal matchd2712d : std_logic := '0';
	
	signal bitvectord2713d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2713d : std_logic := '1';
	signal matchd2713d : std_logic := '0';
	
	signal bitvectord2714d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2714d : std_logic := '0';
	signal matchd2714d : std_logic := '0';
	
	signal bitvectord2715d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2715d : std_logic := '0';
	signal matchd2715d : std_logic := '0';
	
	signal bitvectord2716d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2716d : std_logic := '0';
	signal matchd2716d : std_logic := '0';
	
	signal bitvectord2717d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2717d : std_logic := '0';
	signal matchd2717d : std_logic := '0';
	
	signal bitvectord2718d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2718d : std_logic := '0';
	signal matchd2718d : std_logic := '0';
	
	signal bitvectord2719d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2719d : std_logic := '0';
	signal matchd2719d : std_logic := '0';
	
	signal bitvectord2720d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2720d : std_logic := '0';
	signal matchd2720d : std_logic := '0';
	
	signal bitvectord2721d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2721d : std_logic := '1';
	signal matchd2721d : std_logic := '0';
	
	signal bitvectord2722d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2722d : std_logic := '0';
	signal matchd2722d : std_logic := '0';
	
	signal bitvectord2723d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2723d : std_logic := '0';
	signal matchd2723d : std_logic := '0';
	
	signal bitvectord2724d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2724d : std_logic := '0';
	signal matchd2724d : std_logic := '0';
	
	signal bitvectord2725d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2725d : std_logic := '0';
	signal matchd2725d : std_logic := '0';
	
	signal bitvectord2726d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2726d : std_logic := '0';
	signal matchd2726d : std_logic := '0';
	
	signal bitvectord2727d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2727d : std_logic := '0';
	signal matchd2727d : std_logic := '0';
	
	signal bitvectord2728d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2728d : std_logic := '0';
	signal matchd2728d : std_logic := '0';
	
	signal bitvectord2729d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2729d : std_logic := '0';
	signal matchd2729d : std_logic := '0';
	
	signal bitvectord2730d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2730d : std_logic := '0';
	signal matchd2730d : std_logic := '0';
	
	signal bitvectord2731d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2731d : std_logic := '0';
	signal matchd2731d : std_logic := '0';
	
	signal bitvectord2732d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2732d : std_logic := '0';
	signal matchd2732d : std_logic := '0';
	
	signal bitvectord2733d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2733d : std_logic := '0';
	signal matchd2733d : std_logic := '0';
	
	signal bitvectord2734d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2734d : std_logic := '0';
	signal matchd2734d : std_logic := '0';
	
	signal bitvectord2735d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2735d : std_logic := '0';
	signal matchd2735d : std_logic := '0';
	
	signal bitvectord2736d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2736d : std_logic := '0';
	signal matchd2736d : std_logic := '0';
	
	signal bitvectord2737d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2737d : std_logic := '0';
	signal matchd2737d : std_logic := '0';
	
	signal bitvectord2738d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2738d : std_logic := '0';
	signal matchd2738d : std_logic := '0';
	
	signal bitvectord2739d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2739d : std_logic := '0';
	signal matchd2739d : std_logic := '0';
	
	signal bitvectord2740d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2740d : std_logic := '0';
	signal matchd2740d : std_logic := '0';
	
	signal bitvectord2741d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2741d : std_logic := '0';
	signal matchd2741d : std_logic := '0';
	
	signal bitvectord2742d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2742d : std_logic := '1';
	signal matchd2742d : std_logic := '0';
	
	signal bitvectord2743d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2743d : std_logic := '0';
	signal matchd2743d : std_logic := '0';
	
	signal bitvectord2744d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2744d : std_logic := '0';
	signal matchd2744d : std_logic := '0';
	
	signal bitvectord2745d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2745d : std_logic := '0';
	signal matchd2745d : std_logic := '0';
	
	signal bitvectord2746d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2746d : std_logic := '0';
	signal matchd2746d : std_logic := '0';
	
	signal bitvectord2747d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2747d : std_logic := '0';
	signal matchd2747d : std_logic := '0';
	
	signal bitvectord2748d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2748d : std_logic := '0';
	signal matchd2748d : std_logic := '0';
	
	signal bitvectord2749d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2749d : std_logic := '0';
	signal matchd2749d : std_logic := '0';
	
	signal bitvectord2750d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2750d : std_logic := '0';
	signal matchd2750d : std_logic := '0';
	
	signal bitvectord2751d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2751d : std_logic := '0';
	signal matchd2751d : std_logic := '0';
	
	signal bitvectord2752d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2752d : std_logic := '0';
	signal matchd2752d : std_logic := '0';
	
	signal bitvectord2753d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2753d : std_logic := '0';
	signal matchd2753d : std_logic := '0';
	
	signal bitvectord2754d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2754d : std_logic := '0';
	signal matchd2754d : std_logic := '0';
	
	signal bitvectord2755d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2755d : std_logic := '0';
	signal matchd2755d : std_logic := '0';
	
	signal bitvectord2756d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2756d : std_logic := '0';
	signal matchd2756d : std_logic := '0';
	
	signal bitvectord2757d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2757d : std_logic := '0';
	signal matchd2757d : std_logic := '0';
	
	signal bitvectord2758d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2758d : std_logic := '0';
	signal matchd2758d : std_logic := '0';
	
	signal bitvectord2759d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2759d : std_logic := '0';
	signal matchd2759d : std_logic := '0';
	
	signal bitvectord2760d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2760d : std_logic := '0';
	signal matchd2760d : std_logic := '0';
	
	signal bitvectord2761d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2761d : std_logic := '0';
	signal matchd2761d : std_logic := '0';
	
	signal bitvectord2762d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2762d : std_logic := '0';
	signal matchd2762d : std_logic := '0';
	
	signal bitvectord2763d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2763d : std_logic := '1';
	signal matchd2763d : std_logic := '0';
	
	signal bitvectord2764d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2764d : std_logic := '0';
	signal matchd2764d : std_logic := '0';
	
	signal bitvectord2765d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2765d : std_logic := '0';
	signal matchd2765d : std_logic := '0';
	
	signal bitvectord2766d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2766d : std_logic := '0';
	signal matchd2766d : std_logic := '0';
	
	signal bitvectord2767d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2767d : std_logic := '0';
	signal matchd2767d : std_logic := '0';
	
	signal bitvectord2768d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2768d : std_logic := '0';
	signal matchd2768d : std_logic := '0';
	
	signal bitvectord2769d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2769d : std_logic := '0';
	signal matchd2769d : std_logic := '0';
	
	signal bitvectord2770d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2770d : std_logic := '0';
	signal matchd2770d : std_logic := '0';
	
	signal bitvectord2771d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2771d : std_logic := '0';
	signal matchd2771d : std_logic := '0';
	
	signal bitvectord2772d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2772d : std_logic := '0';
	signal matchd2772d : std_logic := '0';
	
	signal bitvectord2773d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2773d : std_logic := '0';
	signal matchd2773d : std_logic := '0';
	
	signal bitvectord2774d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2774d : std_logic := '0';
	signal matchd2774d : std_logic := '0';
	
	signal bitvectord2775d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2775d : std_logic := '0';
	signal matchd2775d : std_logic := '0';
	
	signal bitvectord2776d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2776d : std_logic := '1';
	signal matchd2776d : std_logic := '0';
	
	signal bitvectord2777d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2777d : std_logic := '0';
	signal matchd2777d : std_logic := '0';
	
	signal bitvectord2778d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2778d : std_logic := '0';
	signal matchd2778d : std_logic := '0';
	
	signal bitvectord2779d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2779d : std_logic := '0';
	signal matchd2779d : std_logic := '0';
	
	signal bitvectord2780d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2780d : std_logic := '0';
	signal matchd2780d : std_logic := '0';
	
	signal bitvectord2781d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2781d : std_logic := '0';
	signal matchd2781d : std_logic := '0';
	
	signal bitvectord2782d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2782d : std_logic := '0';
	signal matchd2782d : std_logic := '0';
	
	signal bitvectord2783d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2783d : std_logic := '0';
	signal matchd2783d : std_logic := '0';
	
	signal bitvectord2784d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2784d : std_logic := '0';
	signal matchd2784d : std_logic := '0';
	
	signal bitvectord2785d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2785d : std_logic := '0';
	signal matchd2785d : std_logic := '0';
	
	signal bitvectord2786d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2786d : std_logic := '0';
	signal matchd2786d : std_logic := '0';
	
	signal bitvectord2787d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2787d : std_logic := '0';
	signal matchd2787d : std_logic := '0';
	
	signal bitvectord2788d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2788d : std_logic := '0';
	signal matchd2788d : std_logic := '0';
	
	signal bitvectord2789d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2789d : std_logic := '0';
	signal matchd2789d : std_logic := '0';
	
	signal bitvectord2790d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2790d : std_logic := '0';
	signal matchd2790d : std_logic := '0';
	
	signal bitvectord2791d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2791d : std_logic := '1';
	signal matchd2791d : std_logic := '0';
	
	signal bitvectord2792d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2792d : std_logic := '0';
	signal matchd2792d : std_logic := '0';
	
	signal bitvectord2793d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2793d : std_logic := '0';
	signal matchd2793d : std_logic := '0';
	
	signal bitvectord2794d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2794d : std_logic := '0';
	signal matchd2794d : std_logic := '0';
	
	signal bitvectord2795d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2795d : std_logic := '0';
	signal matchd2795d : std_logic := '0';
	
	signal bitvectord2796d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2796d : std_logic := '0';
	signal matchd2796d : std_logic := '0';
	
	signal bitvectord2797d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2797d : std_logic := '0';
	signal matchd2797d : std_logic := '0';
	
	signal bitvectord2798d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2798d : std_logic := '0';
	signal matchd2798d : std_logic := '0';
	
	signal bitvectord2799d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2799d : std_logic := '0';
	signal matchd2799d : std_logic := '0';
	
	signal bitvectord2800d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2800d : std_logic := '0';
	signal matchd2800d : std_logic := '0';
	
	signal bitvectord2801d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2801d : std_logic := '0';
	signal matchd2801d : std_logic := '0';
	
	signal bitvectord2802d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2802d : std_logic := '1';
	signal matchd2802d : std_logic := '0';
	
	signal bitvectord2803d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2803d : std_logic := '0';
	signal matchd2803d : std_logic := '0';
	
	signal bitvectord2804d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2804d : std_logic := '0';
	signal matchd2804d : std_logic := '0';
	
	signal bitvectord2805d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2805d : std_logic := '0';
	signal matchd2805d : std_logic := '0';
	
	signal bitvectord2806d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2806d : std_logic := '0';
	signal matchd2806d : std_logic := '0';
	
	signal bitvectord2807d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2807d : std_logic := '0';
	signal matchd2807d : std_logic := '0';
	
	signal bitvectord2808d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2808d : std_logic := '0';
	signal matchd2808d : std_logic := '0';
	
	signal bitvectord2809d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2809d : std_logic := '0';
	signal matchd2809d : std_logic := '0';
	
	signal bitvectord2810d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2810d : std_logic := '0';
	signal matchd2810d : std_logic := '0';
	
	signal bitvectord2811d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2811d : std_logic := '0';
	signal matchd2811d : std_logic := '0';
	
	signal bitvectord2812d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2812d : std_logic := '0';
	signal matchd2812d : std_logic := '0';
	
	signal bitvectord2813d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2813d : std_logic := '0';
	signal matchd2813d : std_logic := '0';
	
	signal bitvectord2814d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2814d : std_logic := '0';
	signal matchd2814d : std_logic := '0';
	
	signal bitvectord2815d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2815d : std_logic := '0';
	signal matchd2815d : std_logic := '0';
	
	signal bitvectord2816d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2816d : std_logic := '0';
	signal matchd2816d : std_logic := '0';
	
	signal bitvectord2817d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2817d : std_logic := '0';
	signal matchd2817d : std_logic := '0';
	
	signal bitvectord2818d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2818d : std_logic := '0';
	signal matchd2818d : std_logic := '0';
	
	signal bitvectord2819d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2819d : std_logic := '1';
	signal matchd2819d : std_logic := '0';
	
	signal bitvectord2820d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2820d : std_logic := '0';
	signal matchd2820d : std_logic := '0';
	
	signal bitvectord2821d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2821d : std_logic := '0';
	signal matchd2821d : std_logic := '0';
	
	signal bitvectord2822d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2822d : std_logic := '0';
	signal matchd2822d : std_logic := '0';
	
	signal bitvectord2823d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2823d : std_logic := '0';
	signal matchd2823d : std_logic := '0';
	
	signal bitvectord2824d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2824d : std_logic := '0';
	signal matchd2824d : std_logic := '0';
	
	signal bitvectord2825d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2825d : std_logic := '0';
	signal matchd2825d : std_logic := '0';
	
	signal bitvectord2826d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2826d : std_logic := '0';
	signal matchd2826d : std_logic := '0';
	
	signal bitvectord2827d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2827d : std_logic := '0';
	signal matchd2827d : std_logic := '0';
	
	signal bitvectord2828d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2828d : std_logic := '0';
	signal matchd2828d : std_logic := '0';
	
	signal bitvectord2829d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2829d : std_logic := '0';
	signal matchd2829d : std_logic := '0';
	
	signal bitvectord2830d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2830d : std_logic := '0';
	signal matchd2830d : std_logic := '0';
	
	signal bitvectord2831d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2831d : std_logic := '0';
	signal matchd2831d : std_logic := '0';
	
	signal bitvectord2832d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2832d : std_logic := '0';
	signal matchd2832d : std_logic := '0';
	
	signal bitvectord2833d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2833d : std_logic := '0';
	signal matchd2833d : std_logic := '0';
	
	signal bitvectord2834d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2834d : std_logic := '0';
	signal matchd2834d : std_logic := '0';
	
	signal bitvectord2835d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2835d : std_logic := '0';
	signal matchd2835d : std_logic := '0';
	
	signal bitvectord2837d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2837d : std_logic := '1';
	signal matchd2837d : std_logic := '0';
	
	signal bitvectord2838d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2838d : std_logic := '0';
	signal matchd2838d : std_logic := '0';
	
	signal bitvectord2839d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2839d : std_logic := '0';
	signal matchd2839d : std_logic := '0';
	
	signal bitvectord2840d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2840d : std_logic := '0';
	signal matchd2840d : std_logic := '0';
	
	signal bitvectord2841d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2841d : std_logic := '0';
	signal matchd2841d : std_logic := '0';
	
	signal bitvectord2842d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2842d : std_logic := '0';
	signal matchd2842d : std_logic := '0';
	
	signal bitvectord2843d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2843d : std_logic := '0';
	signal matchd2843d : std_logic := '0';
	
	signal bitvectord2844d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2844d : std_logic := '0';
	signal matchd2844d : std_logic := '0';
	
	signal bitvectord2845d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2845d : std_logic := '0';
	signal matchd2845d : std_logic := '0';
	
	signal bitvectord2846d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2846d : std_logic := '0';
	signal matchd2846d : std_logic := '0';
	
	signal bitvectord2847d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2847d : std_logic := '0';
	signal matchd2847d : std_logic := '0';
	
	signal bitvectord2848d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2848d : std_logic := '0';
	signal matchd2848d : std_logic := '0';
	
	signal bitvectord2849d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2849d : std_logic := '0';
	signal matchd2849d : std_logic := '0';
	
	signal bitvectord2850d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2850d : std_logic := '0';
	signal matchd2850d : std_logic := '0';
	
	signal bitvectord2851d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2851d : std_logic := '0';
	signal matchd2851d : std_logic := '0';
	
	signal bitvectord2852d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2852d : std_logic := '0';
	signal matchd2852d : std_logic := '0';
	
	signal bitvectord2853d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2853d : std_logic := '1';
	signal matchd2853d : std_logic := '0';
	
	signal bitvectord2854d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2854d : std_logic := '0';
	signal matchd2854d : std_logic := '0';
	
	signal bitvectord2855d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2855d : std_logic := '0';
	signal matchd2855d : std_logic := '0';
	
	signal bitvectord2856d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2856d : std_logic := '0';
	signal matchd2856d : std_logic := '0';
	
	signal bitvectord2857d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2857d : std_logic := '0';
	signal matchd2857d : std_logic := '0';
	
	signal bitvectord2858d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2858d : std_logic := '0';
	signal matchd2858d : std_logic := '0';
	
	signal bitvectord2859d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2859d : std_logic := '0';
	signal matchd2859d : std_logic := '0';
	
	signal bitvectord2860d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2860d : std_logic := '0';
	signal matchd2860d : std_logic := '0';
	
	signal bitvectord2861d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled2861d : std_logic := '0';
	signal matchd2861d : std_logic := '0';
	
	signal bitvectord2862d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2862d : std_logic := '0';
	signal matchd2862d : std_logic := '0';
	
	signal bitvectord2863d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2863d : std_logic := '0';
	signal matchd2863d : std_logic := '0';
	
	signal bitvectord2864d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2864d : std_logic := '0';
	signal matchd2864d : std_logic := '0';
	
	signal bitvectord2865d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2865d : std_logic := '0';
	signal matchd2865d : std_logic := '0';
	
	signal bitvectord2866d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2866d : std_logic := '0';
	signal matchd2866d : std_logic := '0';
	
	signal bitvectord2867d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2867d : std_logic := '0';
	signal matchd2867d : std_logic := '0';
	
	signal bitvectord2868d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2868d : std_logic := '0';
	signal matchd2868d : std_logic := '0';
	
	signal bitvectord2870d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2870d : std_logic := '1';
	signal matchd2870d : std_logic := '0';
	
	signal bitvectord2871d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2871d : std_logic := '0';
	signal matchd2871d : std_logic := '0';
	
	signal bitvectord2872d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2872d : std_logic := '0';
	signal matchd2872d : std_logic := '0';
	
	signal bitvectord2873d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2873d : std_logic := '0';
	signal matchd2873d : std_logic := '0';
	
	signal bitvectord2874d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2874d : std_logic := '0';
	signal matchd2874d : std_logic := '0';
	
	signal bitvectord2875d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2875d : std_logic := '0';
	signal matchd2875d : std_logic := '0';
	
	signal bitvectord2876d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2876d : std_logic := '0';
	signal matchd2876d : std_logic := '0';
	
	signal bitvectord2877d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2877d : std_logic := '0';
	signal matchd2877d : std_logic := '0';
	
	signal bitvectord2878d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2878d : std_logic := '0';
	signal matchd2878d : std_logic := '0';
	
	signal bitvectord2879d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2879d : std_logic := '0';
	signal matchd2879d : std_logic := '0';
	
	signal bitvectord2880d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2880d : std_logic := '0';
	signal matchd2880d : std_logic := '0';
	
	signal bitvectord2881d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2881d : std_logic := '0';
	signal matchd2881d : std_logic := '0';
	
	signal bitvectord2882d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2882d : std_logic := '0';
	signal matchd2882d : std_logic := '0';
	
	signal bitvectord2883d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2883d : std_logic := '1';
	signal matchd2883d : std_logic := '0';
	
	signal bitvectord2884d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2884d : std_logic := '0';
	signal matchd2884d : std_logic := '0';
	
	signal bitvectord2885d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2885d : std_logic := '0';
	signal matchd2885d : std_logic := '0';
	
	signal bitvectord2886d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2886d : std_logic := '0';
	signal matchd2886d : std_logic := '0';
	
	signal bitvectord2887d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2887d : std_logic := '0';
	signal matchd2887d : std_logic := '0';
	
	signal bitvectord2888d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2888d : std_logic := '0';
	signal matchd2888d : std_logic := '0';
	
	signal bitvectord2889d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2889d : std_logic := '0';
	signal matchd2889d : std_logic := '0';
	
	signal bitvectord2890d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2890d : std_logic := '0';
	signal matchd2890d : std_logic := '0';
	
	signal bitvectord2891d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2891d : std_logic := '0';
	signal matchd2891d : std_logic := '0';
	
	signal bitvectord2892d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2892d : std_logic := '0';
	signal matchd2892d : std_logic := '0';
	
	signal bitvectord2893d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2893d : std_logic := '0';
	signal matchd2893d : std_logic := '0';
	
	signal bitvectord2894d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2894d : std_logic := '0';
	signal matchd2894d : std_logic := '0';
	
	signal bitvectord2895d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2895d : std_logic := '0';
	signal matchd2895d : std_logic := '0';
	
	signal bitvectord2896d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2896d : std_logic := '0';
	signal matchd2896d : std_logic := '0';
	
	signal bitvectord2897d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2897d : std_logic := '0';
	signal matchd2897d : std_logic := '0';
	
	signal bitvectord2898d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2898d : std_logic := '0';
	signal matchd2898d : std_logic := '0';
	
	signal bitvectord2899d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2899d : std_logic := '0';
	signal matchd2899d : std_logic := '0';
	
	signal bitvectord2900d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2900d : std_logic := '1';
	signal matchd2900d : std_logic := '0';
	
	signal bitvectord2901d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2901d : std_logic := '0';
	signal matchd2901d : std_logic := '0';
	
	signal bitvectord2902d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2902d : std_logic := '0';
	signal matchd2902d : std_logic := '0';
	
	signal bitvectord2903d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2903d : std_logic := '0';
	signal matchd2903d : std_logic := '0';
	
	signal bitvectord2904d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2904d : std_logic := '0';
	signal matchd2904d : std_logic := '0';
	
	signal bitvectord2905d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2905d : std_logic := '0';
	signal matchd2905d : std_logic := '0';
	
	signal bitvectord2906d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2906d : std_logic := '0';
	signal matchd2906d : std_logic := '0';
	
	signal bitvectord2907d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2907d : std_logic := '0';
	signal matchd2907d : std_logic := '0';
	
	signal bitvectord2908d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2908d : std_logic := '0';
	signal matchd2908d : std_logic := '0';
	
	signal bitvectord2909d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2909d : std_logic := '0';
	signal matchd2909d : std_logic := '0';
	
	signal bitvectord2910d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2910d : std_logic := '0';
	signal matchd2910d : std_logic := '0';
	
	signal bitvectord2911d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2911d : std_logic := '0';
	signal matchd2911d : std_logic := '0';
	
	signal bitvectord2912d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2912d : std_logic := '0';
	signal matchd2912d : std_logic := '0';
	
	signal bitvectord2913d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2913d : std_logic := '1';
	signal matchd2913d : std_logic := '0';
	
	signal bitvectord2914d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2914d : std_logic := '0';
	signal matchd2914d : std_logic := '0';
	
	signal bitvectord2915d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2915d : std_logic := '0';
	signal matchd2915d : std_logic := '0';
	
	signal bitvectord2916d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2916d : std_logic := '0';
	signal matchd2916d : std_logic := '0';
	
	signal bitvectord2917d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2917d : std_logic := '0';
	signal matchd2917d : std_logic := '0';
	
	signal bitvectord2918d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2918d : std_logic := '0';
	signal matchd2918d : std_logic := '0';
	
	signal bitvectord2919d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2919d : std_logic := '0';
	signal matchd2919d : std_logic := '0';
	
	signal bitvectord2920d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2920d : std_logic := '0';
	signal matchd2920d : std_logic := '0';
	
	signal bitvectord2921d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2921d : std_logic := '0';
	signal matchd2921d : std_logic := '0';
	
	signal bitvectord2922d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2922d : std_logic := '0';
	signal matchd2922d : std_logic := '0';
	
	signal bitvectord2923d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2923d : std_logic := '0';
	signal matchd2923d : std_logic := '0';
	
	signal bitvectord2924d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2924d : std_logic := '0';
	signal matchd2924d : std_logic := '0';
	
	signal bitvectord2925d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2925d : std_logic := '1';
	signal matchd2925d : std_logic := '0';
	
	signal bitvectord2926d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2926d : std_logic := '0';
	signal matchd2926d : std_logic := '0';
	
	signal bitvectord2927d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2927d : std_logic := '0';
	signal matchd2927d : std_logic := '0';
	
	signal bitvectord2928d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2928d : std_logic := '0';
	signal matchd2928d : std_logic := '0';
	
	signal bitvectord2929d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2929d : std_logic := '0';
	signal matchd2929d : std_logic := '0';
	
	signal bitvectord2930d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2930d : std_logic := '0';
	signal matchd2930d : std_logic := '0';
	
	signal bitvectord2931d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2931d : std_logic := '0';
	signal matchd2931d : std_logic := '0';
	
	signal bitvectord2932d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2932d : std_logic := '0';
	signal matchd2932d : std_logic := '0';
	
	signal bitvectord2933d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2933d : std_logic := '0';
	signal matchd2933d : std_logic := '0';
	
	signal bitvectord2934d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2934d : std_logic := '0';
	signal matchd2934d : std_logic := '0';
	
	signal bitvectord2935d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2935d : std_logic := '0';
	signal matchd2935d : std_logic := '0';
	
	signal bitvectord2936d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2936d : std_logic := '0';
	signal matchd2936d : std_logic := '0';
	
	signal bitvectord2937d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2937d : std_logic := '0';
	signal matchd2937d : std_logic := '0';
	
	signal bitvectord2938d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2938d : std_logic := '0';
	signal matchd2938d : std_logic := '0';
	
	signal bitvectord2939d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2939d : std_logic := '0';
	signal matchd2939d : std_logic := '0';
	
	signal bitvectord2940d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2940d : std_logic := '0';
	signal matchd2940d : std_logic := '0';
	
	signal bitvectord2941d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2941d : std_logic := '0';
	signal matchd2941d : std_logic := '0';
	
	signal bitvectord2942d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2942d : std_logic := '1';
	signal matchd2942d : std_logic := '0';
	
	signal bitvectord2943d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2943d : std_logic := '0';
	signal matchd2943d : std_logic := '0';
	
	signal bitvectord2944d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2944d : std_logic := '0';
	signal matchd2944d : std_logic := '0';
	
	signal bitvectord2945d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2945d : std_logic := '0';
	signal matchd2945d : std_logic := '0';
	
	signal bitvectord2946d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2946d : std_logic := '0';
	signal matchd2946d : std_logic := '0';
	
	signal bitvectord2947d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2947d : std_logic := '0';
	signal matchd2947d : std_logic := '0';
	
	signal bitvectord2948d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2948d : std_logic := '0';
	signal matchd2948d : std_logic := '0';
	
	signal bitvectord2949d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2949d : std_logic := '0';
	signal matchd2949d : std_logic := '0';
	
	signal bitvectord2950d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2950d : std_logic := '0';
	signal matchd2950d : std_logic := '0';
	
	signal bitvectord2951d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2951d : std_logic := '0';
	signal matchd2951d : std_logic := '0';
	
	signal bitvectord2952d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2952d : std_logic := '0';
	signal matchd2952d : std_logic := '0';
	
	signal bitvectord2953d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2953d : std_logic := '0';
	signal matchd2953d : std_logic := '0';
	
	signal bitvectord2954d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2954d : std_logic := '0';
	signal matchd2954d : std_logic := '0';
	
	signal bitvectord2955d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2955d : std_logic := '0';
	signal matchd2955d : std_logic := '0';
	
	signal bitvectord2956d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2956d : std_logic := '0';
	signal matchd2956d : std_logic := '0';
	
	signal bitvectord2957d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2957d : std_logic := '1';
	signal matchd2957d : std_logic := '0';
	
	signal bitvectord2958d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2958d : std_logic := '0';
	signal matchd2958d : std_logic := '0';
	
	signal bitvectord2959d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2959d : std_logic := '0';
	signal matchd2959d : std_logic := '0';
	
	signal bitvectord2960d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2960d : std_logic := '0';
	signal matchd2960d : std_logic := '0';
	
	signal bitvectord2961d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2961d : std_logic := '0';
	signal matchd2961d : std_logic := '0';
	
	signal bitvectord2962d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2962d : std_logic := '0';
	signal matchd2962d : std_logic := '0';
	
	signal bitvectord2963d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2963d : std_logic := '0';
	signal matchd2963d : std_logic := '0';
	
	signal bitvectord2964d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2964d : std_logic := '0';
	signal matchd2964d : std_logic := '0';
	
	signal bitvectord2965d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2965d : std_logic := '0';
	signal matchd2965d : std_logic := '0';
	
	signal bitvectord2966d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2966d : std_logic := '0';
	signal matchd2966d : std_logic := '0';
	
	signal bitvectord2967d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2967d : std_logic := '0';
	signal matchd2967d : std_logic := '0';
	
	signal bitvectord2968d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2968d : std_logic := '1';
	signal matchd2968d : std_logic := '0';
	
	signal bitvectord2969d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2969d : std_logic := '0';
	signal matchd2969d : std_logic := '0';
	
	signal bitvectord2970d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2970d : std_logic := '0';
	signal matchd2970d : std_logic := '0';
	
	signal bitvectord2971d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2971d : std_logic := '0';
	signal matchd2971d : std_logic := '0';
	
	signal bitvectord2972d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2972d : std_logic := '0';
	signal matchd2972d : std_logic := '0';
	
	signal bitvectord2973d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2973d : std_logic := '0';
	signal matchd2973d : std_logic := '0';
	
	signal bitvectord2974d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2974d : std_logic := '0';
	signal matchd2974d : std_logic := '0';
	
	signal bitvectord2975d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2975d : std_logic := '0';
	signal matchd2975d : std_logic := '0';
	
	signal bitvectord2976d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2976d : std_logic := '0';
	signal matchd2976d : std_logic := '0';
	
	signal bitvectord2977d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2977d : std_logic := '0';
	signal matchd2977d : std_logic := '0';
	
	signal bitvectord2978d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2978d : std_logic := '0';
	signal matchd2978d : std_logic := '0';
	
	signal bitvectord2979d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2979d : std_logic := '0';
	signal matchd2979d : std_logic := '0';
	
	signal bitvectord2980d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2980d : std_logic := '1';
	signal matchd2980d : std_logic := '0';
	
	signal bitvectord2981d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2981d : std_logic := '0';
	signal matchd2981d : std_logic := '0';
	
	signal bitvectord2982d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2982d : std_logic := '0';
	signal matchd2982d : std_logic := '0';
	
	signal bitvectord2983d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2983d : std_logic := '0';
	signal matchd2983d : std_logic := '0';
	
	signal bitvectord2984d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2984d : std_logic := '0';
	signal matchd2984d : std_logic := '0';
	
	signal bitvectord2985d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2985d : std_logic := '0';
	signal matchd2985d : std_logic := '0';
	
	signal bitvectord2986d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000";
	signal Enabled2986d : std_logic := '0';
	signal matchd2986d : std_logic := '0';
	
	signal bitvectord2987d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2987d : std_logic := '0';
	signal matchd2987d : std_logic := '0';
	
	signal bitvectord2988d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled2988d : std_logic := '0';
	signal matchd2988d : std_logic := '0';
	
	signal bitvectord2989d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2989d : std_logic := '0';
	signal matchd2989d : std_logic := '0';
	
	signal bitvectord2990d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2990d : std_logic := '0';
	signal matchd2990d : std_logic := '0';
	
	signal bitvectord2991d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2991d : std_logic := '0';
	signal matchd2991d : std_logic := '0';
	
	signal bitvectord2992d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2992d : std_logic := '0';
	signal matchd2992d : std_logic := '0';
	
	signal bitvectord2993d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2993d : std_logic := '0';
	signal matchd2993d : std_logic := '0';
	
	signal bitvectord2994d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled2994d : std_logic := '1';
	signal matchd2994d : std_logic := '0';
	
	signal bitvectord2995d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2995d : std_logic := '0';
	signal matchd2995d : std_logic := '0';
	
	signal bitvectord2996d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2996d : std_logic := '0';
	signal matchd2996d : std_logic := '0';
	
	signal bitvectord2997d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2997d : std_logic := '0';
	signal matchd2997d : std_logic := '0';
	
	signal bitvectord2998d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled2998d : std_logic := '0';
	signal matchd2998d : std_logic := '0';
	
	signal bitvectord2999d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled2999d : std_logic := '0';
	signal matchd2999d : std_logic := '0';
	
	signal bitvectord3000d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3000d : std_logic := '0';
	signal matchd3000d : std_logic := '0';
	
	signal bitvectord3001d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3001d : std_logic := '0';
	signal matchd3001d : std_logic := '0';
	
	signal bitvectord3002d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3002d : std_logic := '0';
	signal matchd3002d : std_logic := '0';
	
	signal bitvectord3003d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3003d : std_logic := '0';
	signal matchd3003d : std_logic := '0';
	
	signal bitvectord3004d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3004d : std_logic := '0';
	signal matchd3004d : std_logic := '0';
	
	signal bitvectord3005d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3005d : std_logic := '0';
	signal matchd3005d : std_logic := '0';
	
	signal bitvectord3006d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3006d : std_logic := '0';
	signal matchd3006d : std_logic := '0';
	
	signal bitvectord3007d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3007d : std_logic := '0';
	signal matchd3007d : std_logic := '0';
	
	signal bitvectord3008d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3008d : std_logic := '1';
	signal matchd3008d : std_logic := '0';
	
	signal bitvectord3009d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3009d : std_logic := '0';
	signal matchd3009d : std_logic := '0';
	
	signal bitvectord3010d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3010d : std_logic := '0';
	signal matchd3010d : std_logic := '0';
	
	signal bitvectord3011d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3011d : std_logic := '0';
	signal matchd3011d : std_logic := '0';
	
	signal bitvectord3012d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3012d : std_logic := '0';
	signal matchd3012d : std_logic := '0';
	
	signal bitvectord3013d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3013d : std_logic := '0';
	signal matchd3013d : std_logic := '0';
	
	signal bitvectord3014d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000";
	signal Enabled3014d : std_logic := '0';
	signal matchd3014d : std_logic := '0';
	
	signal bitvectord3015d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3015d : std_logic := '0';
	signal matchd3015d : std_logic := '0';
	
	signal bitvectord3016d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3016d : std_logic := '0';
	signal matchd3016d : std_logic := '0';
	
	signal bitvectord3017d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3017d : std_logic := '0';
	signal matchd3017d : std_logic := '0';
	
	signal bitvectord3018d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3018d : std_logic := '0';
	signal matchd3018d : std_logic := '0';
	
	signal bitvectord3019d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3019d : std_logic := '0';
	signal matchd3019d : std_logic := '0';
	
	signal bitvectord3020d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3020d : std_logic := '0';
	signal matchd3020d : std_logic := '0';
	
	signal bitvectord3021d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3021d : std_logic := '0';
	signal matchd3021d : std_logic := '0';
	
	signal bitvectord3022d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3022d : std_logic := '0';
	signal matchd3022d : std_logic := '0';
	
	signal bitvectord3023d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3023d : std_logic := '0';
	signal matchd3023d : std_logic := '0';
	
	signal bitvectord3024d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3024d : std_logic := '1';
	signal matchd3024d : std_logic := '0';
	
	signal bitvectord3025d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3025d : std_logic := '0';
	signal matchd3025d : std_logic := '0';
	
	signal bitvectord3026d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3026d : std_logic := '0';
	signal matchd3026d : std_logic := '0';
	
	signal bitvectord3027d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3027d : std_logic := '0';
	signal matchd3027d : std_logic := '0';
	
	signal bitvectord3028d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3028d : std_logic := '0';
	signal matchd3028d : std_logic := '0';
	
	signal bitvectord3029d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3029d : std_logic := '0';
	signal matchd3029d : std_logic := '0';
	
	signal bitvectord3030d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3030d : std_logic := '0';
	signal matchd3030d : std_logic := '0';
	
	signal bitvectord3031d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3031d : std_logic := '0';
	signal matchd3031d : std_logic := '0';
	
	signal bitvectord3032d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3032d : std_logic := '0';
	signal matchd3032d : std_logic := '0';
	
	signal bitvectord3033d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3033d : std_logic := '0';
	signal matchd3033d : std_logic := '0';
	
	signal bitvectord3034d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3034d : std_logic := '0';
	signal matchd3034d : std_logic := '0';
	
	signal bitvectord3035d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3035d : std_logic := '0';
	signal matchd3035d : std_logic := '0';
	
	signal bitvectord3036d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3036d : std_logic := '0';
	signal matchd3036d : std_logic := '0';
	
	signal bitvectord3037d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3037d : std_logic := '0';
	signal matchd3037d : std_logic := '0';
	
	signal bitvectord3038d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3038d : std_logic := '0';
	signal matchd3038d : std_logic := '0';
	
	signal bitvectord3039d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3039d : std_logic := '0';
	signal matchd3039d : std_logic := '0';
	
	signal bitvectord3040d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3040d : std_logic := '0';
	signal matchd3040d : std_logic := '0';
	
	signal bitvectord3041d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3041d : std_logic := '1';
	signal matchd3041d : std_logic := '0';
	
	signal bitvectord3042d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3042d : std_logic := '0';
	signal matchd3042d : std_logic := '0';
	
	signal bitvectord3043d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3043d : std_logic := '0';
	signal matchd3043d : std_logic := '0';
	
	signal bitvectord3044d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3044d : std_logic := '0';
	signal matchd3044d : std_logic := '0';
	
	signal bitvectord3045d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3045d : std_logic := '0';
	signal matchd3045d : std_logic := '0';
	
	signal bitvectord3046d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3046d : std_logic := '0';
	signal matchd3046d : std_logic := '0';
	
	signal bitvectord3047d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3047d : std_logic := '0';
	signal matchd3047d : std_logic := '0';
	
	signal bitvectord3048d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3048d : std_logic := '0';
	signal matchd3048d : std_logic := '0';
	
	signal bitvectord3049d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3049d : std_logic := '0';
	signal matchd3049d : std_logic := '0';
	
	signal bitvectord3050d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3050d : std_logic := '0';
	signal matchd3050d : std_logic := '0';
	
	signal bitvectord3051d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3051d : std_logic := '0';
	signal matchd3051d : std_logic := '0';
	
	signal bitvectord3052d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3052d : std_logic := '0';
	signal matchd3052d : std_logic := '0';
	
	signal bitvectord3053d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3053d : std_logic := '0';
	signal matchd3053d : std_logic := '0';
	
	signal bitvectord3054d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3054d : std_logic := '0';
	signal matchd3054d : std_logic := '0';
	
	signal bitvectord3055d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3055d : std_logic := '0';
	signal matchd3055d : std_logic := '0';
	
	signal bitvectord3056d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3056d : std_logic := '0';
	signal matchd3056d : std_logic := '0';
	
	signal bitvectord3057d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3057d : std_logic := '0';
	signal matchd3057d : std_logic := '0';
	
	signal bitvectord3059d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3059d : std_logic := '1';
	signal matchd3059d : std_logic := '0';
	
	signal bitvectord3060d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3060d : std_logic := '0';
	signal matchd3060d : std_logic := '0';
	
	signal bitvectord3061d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3061d : std_logic := '0';
	signal matchd3061d : std_logic := '0';
	
	signal bitvectord3062d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3062d : std_logic := '0';
	signal matchd3062d : std_logic := '0';
	
	signal bitvectord3063d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3063d : std_logic := '0';
	signal matchd3063d : std_logic := '0';
	
	signal bitvectord3064d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3064d : std_logic := '0';
	signal matchd3064d : std_logic := '0';
	
	signal bitvectord3065d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3065d : std_logic := '0';
	signal matchd3065d : std_logic := '0';
	
	signal bitvectord3066d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3066d : std_logic := '0';
	signal matchd3066d : std_logic := '0';
	
	signal bitvectord3067d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3067d : std_logic := '0';
	signal matchd3067d : std_logic := '0';
	
	signal bitvectord3068d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3068d : std_logic := '0';
	signal matchd3068d : std_logic := '0';
	
	signal bitvectord3069d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3069d : std_logic := '0';
	signal matchd3069d : std_logic := '0';
	
	signal bitvectord3070d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3070d : std_logic := '0';
	signal matchd3070d : std_logic := '0';
	
	signal bitvectord3071d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3071d : std_logic := '0';
	signal matchd3071d : std_logic := '0';
	
	signal bitvectord3072d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3072d : std_logic := '0';
	signal matchd3072d : std_logic := '0';
	
	signal bitvectord3073d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3073d : std_logic := '0';
	signal matchd3073d : std_logic := '0';
	
	signal bitvectord3074d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3074d : std_logic := '0';
	signal matchd3074d : std_logic := '0';
	
	signal bitvectord3075d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3075d : std_logic := '0';
	signal matchd3075d : std_logic := '0';
	
	signal bitvectord3076d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3076d : std_logic := '0';
	signal matchd3076d : std_logic := '0';
	
	signal bitvectord3077d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3077d : std_logic := '0';
	signal matchd3077d : std_logic := '0';
	
	signal bitvectord3078d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3078d : std_logic := '1';
	signal matchd3078d : std_logic := '0';
	
	signal bitvectord3079d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3079d : std_logic := '0';
	signal matchd3079d : std_logic := '0';
	
	signal bitvectord3080d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3080d : std_logic := '0';
	signal matchd3080d : std_logic := '0';
	
	signal bitvectord3081d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3081d : std_logic := '0';
	signal matchd3081d : std_logic := '0';
	
	signal bitvectord3082d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3082d : std_logic := '0';
	signal matchd3082d : std_logic := '0';
	
	signal bitvectord3083d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3083d : std_logic := '0';
	signal matchd3083d : std_logic := '0';
	
	signal bitvectord3084d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3084d : std_logic := '0';
	signal matchd3084d : std_logic := '0';
	
	signal bitvectord3085d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3085d : std_logic := '0';
	signal matchd3085d : std_logic := '0';
	
	signal bitvectord3086d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3086d : std_logic := '0';
	signal matchd3086d : std_logic := '0';
	
	signal bitvectord3087d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3087d : std_logic := '0';
	signal matchd3087d : std_logic := '0';
	
	signal bitvectord3088d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3088d : std_logic := '0';
	signal matchd3088d : std_logic := '0';
	
	signal bitvectord3089d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3089d : std_logic := '0';
	signal matchd3089d : std_logic := '0';
	
	signal bitvectord3090d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3090d : std_logic := '0';
	signal matchd3090d : std_logic := '0';
	
	signal bitvectord3091d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3091d : std_logic := '0';
	signal matchd3091d : std_logic := '0';
	
	signal bitvectord3092d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3092d : std_logic := '0';
	signal matchd3092d : std_logic := '0';
	
	signal bitvectord3093d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3093d : std_logic := '0';
	signal matchd3093d : std_logic := '0';
	
	signal bitvectord3094d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3094d : std_logic := '0';
	signal matchd3094d : std_logic := '0';
	
	signal bitvectord3095d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3095d : std_logic := '0';
	signal matchd3095d : std_logic := '0';
	
	signal bitvectord3096d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3096d : std_logic := '0';
	signal matchd3096d : std_logic := '0';
	
	signal bitvectord3097d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3097d : std_logic := '1';
	signal matchd3097d : std_logic := '0';
	
	signal bitvectord3098d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3098d : std_logic := '0';
	signal matchd3098d : std_logic := '0';
	
	signal bitvectord3099d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3099d : std_logic := '0';
	signal matchd3099d : std_logic := '0';
	
	signal bitvectord3100d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3100d : std_logic := '0';
	signal matchd3100d : std_logic := '0';
	
	signal bitvectord3101d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3101d : std_logic := '0';
	signal matchd3101d : std_logic := '0';
	
	signal bitvectord3102d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3102d : std_logic := '0';
	signal matchd3102d : std_logic := '0';
	
	signal bitvectord3103d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3103d : std_logic := '0';
	signal matchd3103d : std_logic := '0';
	
	signal bitvectord3104d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3104d : std_logic := '0';
	signal matchd3104d : std_logic := '0';
	
	signal bitvectord3105d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3105d : std_logic := '0';
	signal matchd3105d : std_logic := '0';
	
	signal bitvectord3106d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3106d : std_logic := '0';
	signal matchd3106d : std_logic := '0';
	
	signal bitvectord3107d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3107d : std_logic := '0';
	signal matchd3107d : std_logic := '0';
	
	signal bitvectord3108d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3108d : std_logic := '0';
	signal matchd3108d : std_logic := '0';
	
	signal bitvectord3109d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3109d : std_logic := '0';
	signal matchd3109d : std_logic := '0';
	
	signal bitvectord3110d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3110d : std_logic := '0';
	signal matchd3110d : std_logic := '0';
	
	signal bitvectord3111d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3111d : std_logic := '0';
	signal matchd3111d : std_logic := '0';
	
	signal bitvectord3112d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3112d : std_logic := '0';
	signal matchd3112d : std_logic := '0';
	
	signal bitvectord3113d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3113d : std_logic := '0';
	signal matchd3113d : std_logic := '0';
	
	signal bitvectord3114d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3114d : std_logic := '0';
	signal matchd3114d : std_logic := '0';
	
	signal bitvectord3115d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3115d : std_logic := '0';
	signal matchd3115d : std_logic := '0';
	
	signal bitvectord3117d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3117d : std_logic := '1';
	signal matchd3117d : std_logic := '0';
	
	signal bitvectord3118d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3118d : std_logic := '0';
	signal matchd3118d : std_logic := '0';
	
	signal bitvectord3119d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3119d : std_logic := '0';
	signal matchd3119d : std_logic := '0';
	
	signal bitvectord3120d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3120d : std_logic := '0';
	signal matchd3120d : std_logic := '0';
	
	signal bitvectord3121d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3121d : std_logic := '0';
	signal matchd3121d : std_logic := '0';
	
	signal bitvectord3122d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3122d : std_logic := '0';
	signal matchd3122d : std_logic := '0';
	
	signal bitvectord3123d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000";
	signal Enabled3123d : std_logic := '0';
	signal matchd3123d : std_logic := '0';
	
	signal bitvectord3124d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3124d : std_logic := '0';
	signal matchd3124d : std_logic := '0';
	
	signal bitvectord3125d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3125d : std_logic := '0';
	signal matchd3125d : std_logic := '0';
	
	signal bitvectord3126d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3126d : std_logic := '0';
	signal matchd3126d : std_logic := '0';
	
	signal bitvectord3127d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3127d : std_logic := '0';
	signal matchd3127d : std_logic := '0';
	
	signal bitvectord3128d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3128d : std_logic := '0';
	signal matchd3128d : std_logic := '0';
	
	signal bitvectord3129d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3129d : std_logic := '0';
	signal matchd3129d : std_logic := '0';
	
	signal bitvectord3130d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3130d : std_logic := '0';
	signal matchd3130d : std_logic := '0';
	
	signal bitvectord3131d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3131d : std_logic := '1';
	signal matchd3131d : std_logic := '0';
	
	signal bitvectord3132d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3132d : std_logic := '0';
	signal matchd3132d : std_logic := '0';
	
	signal bitvectord3133d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3133d : std_logic := '0';
	signal matchd3133d : std_logic := '0';
	
	signal bitvectord3134d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3134d : std_logic := '0';
	signal matchd3134d : std_logic := '0';
	
	signal bitvectord3135d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3135d : std_logic := '0';
	signal matchd3135d : std_logic := '0';
	
	signal bitvectord3136d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3136d : std_logic := '0';
	signal matchd3136d : std_logic := '0';
	
	signal bitvectord3137d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3137d : std_logic := '0';
	signal matchd3137d : std_logic := '0';
	
	signal bitvectord3138d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3138d : std_logic := '0';
	signal matchd3138d : std_logic := '0';
	
	signal bitvectord3139d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3139d : std_logic := '0';
	signal matchd3139d : std_logic := '0';
	
	signal bitvectord3140d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3140d : std_logic := '0';
	signal matchd3140d : std_logic := '0';
	
	signal bitvectord3141d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3141d : std_logic := '0';
	signal matchd3141d : std_logic := '0';
	
	signal bitvectord3142d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3142d : std_logic := '0';
	signal matchd3142d : std_logic := '0';
	
	signal bitvectord3143d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3143d : std_logic := '0';
	signal matchd3143d : std_logic := '0';
	
	signal bitvectord3144d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3144d : std_logic := '0';
	signal matchd3144d : std_logic := '0';
	
	signal bitvectord3145d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3145d : std_logic := '0';
	signal matchd3145d : std_logic := '0';
	
	signal bitvectord3146d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3146d : std_logic := '0';
	signal matchd3146d : std_logic := '0';
	
	signal bitvectord3147d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3147d : std_logic := '0';
	signal matchd3147d : std_logic := '0';
	
	signal bitvectord3148d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3148d : std_logic := '0';
	signal matchd3148d : std_logic := '0';
	
	signal bitvectord3149d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3149d : std_logic := '0';
	signal matchd3149d : std_logic := '0';
	
	signal bitvectord3150d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3150d : std_logic := '1';
	signal matchd3150d : std_logic := '0';
	
	signal bitvectord3151d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3151d : std_logic := '0';
	signal matchd3151d : std_logic := '0';
	
	signal bitvectord3152d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3152d : std_logic := '0';
	signal matchd3152d : std_logic := '0';
	
	signal bitvectord3153d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3153d : std_logic := '0';
	signal matchd3153d : std_logic := '0';
	
	signal bitvectord3154d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3154d : std_logic := '0';
	signal matchd3154d : std_logic := '0';
	
	signal bitvectord3155d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3155d : std_logic := '0';
	signal matchd3155d : std_logic := '0';
	
	signal bitvectord3156d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3156d : std_logic := '0';
	signal matchd3156d : std_logic := '0';
	
	signal bitvectord3157d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3157d : std_logic := '0';
	signal matchd3157d : std_logic := '0';
	
	signal bitvectord3158d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3158d : std_logic := '0';
	signal matchd3158d : std_logic := '0';
	
	signal bitvectord3159d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3159d : std_logic := '0';
	signal matchd3159d : std_logic := '0';
	
	signal bitvectord3160d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3160d : std_logic := '0';
	signal matchd3160d : std_logic := '0';
	
	signal bitvectord3161d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3161d : std_logic := '0';
	signal matchd3161d : std_logic := '0';
	
	signal bitvectord3162d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3162d : std_logic := '0';
	signal matchd3162d : std_logic := '0';
	
	signal bitvectord3163d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3163d : std_logic := '0';
	signal matchd3163d : std_logic := '0';
	
	signal bitvectord3164d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3164d : std_logic := '0';
	signal matchd3164d : std_logic := '0';
	
	signal bitvectord3165d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3165d : std_logic := '0';
	signal matchd3165d : std_logic := '0';
	
	signal bitvectord3166d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3166d : std_logic := '1';
	signal matchd3166d : std_logic := '0';
	
	signal bitvectord3167d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3167d : std_logic := '0';
	signal matchd3167d : std_logic := '0';
	
	signal bitvectord3168d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3168d : std_logic := '0';
	signal matchd3168d : std_logic := '0';
	
	signal bitvectord3169d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3169d : std_logic := '0';
	signal matchd3169d : std_logic := '0';
	
	signal bitvectord3170d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3170d : std_logic := '0';
	signal matchd3170d : std_logic := '0';
	
	signal bitvectord3171d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3171d : std_logic := '0';
	signal matchd3171d : std_logic := '0';
	
	signal bitvectord3172d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3172d : std_logic := '0';
	signal matchd3172d : std_logic := '0';
	
	signal bitvectord3173d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3173d : std_logic := '0';
	signal matchd3173d : std_logic := '0';
	
	signal bitvectord3174d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3174d : std_logic := '0';
	signal matchd3174d : std_logic := '0';
	
	signal bitvectord3175d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3175d : std_logic := '0';
	signal matchd3175d : std_logic := '0';
	
	signal bitvectord3176d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3176d : std_logic := '0';
	signal matchd3176d : std_logic := '0';
	
	signal bitvectord3177d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3177d : std_logic := '0';
	signal matchd3177d : std_logic := '0';
	
	signal bitvectord3178d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3178d : std_logic := '0';
	signal matchd3178d : std_logic := '0';
	
	signal bitvectord3179d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3179d : std_logic := '0';
	signal matchd3179d : std_logic := '0';
	
	signal bitvectord3180d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3180d : std_logic := '0';
	signal matchd3180d : std_logic := '0';
	
	signal bitvectord3181d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3181d : std_logic := '0';
	signal matchd3181d : std_logic := '0';
	
	signal bitvectord3183d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3183d : std_logic := '1';
	signal matchd3183d : std_logic := '0';
	
	signal bitvectord3184d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3184d : std_logic := '0';
	signal matchd3184d : std_logic := '0';
	
	signal bitvectord3185d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3185d : std_logic := '0';
	signal matchd3185d : std_logic := '0';
	
	signal bitvectord3186d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3186d : std_logic := '0';
	signal matchd3186d : std_logic := '0';
	
	signal bitvectord3187d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3187d : std_logic := '0';
	signal matchd3187d : std_logic := '0';
	
	signal bitvectord3188d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3188d : std_logic := '0';
	signal matchd3188d : std_logic := '0';
	
	signal bitvectord3189d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3189d : std_logic := '0';
	signal matchd3189d : std_logic := '0';
	
	signal bitvectord3190d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3190d : std_logic := '0';
	signal matchd3190d : std_logic := '0';
	
	signal bitvectord3191d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3191d : std_logic := '0';
	signal matchd3191d : std_logic := '0';
	
	signal bitvectord3192d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3192d : std_logic := '0';
	signal matchd3192d : std_logic := '0';
	
	signal bitvectord3193d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3193d : std_logic := '0';
	signal matchd3193d : std_logic := '0';
	
	signal bitvectord3194d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3194d : std_logic := '0';
	signal matchd3194d : std_logic := '0';
	
	signal bitvectord3195d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3195d : std_logic := '0';
	signal matchd3195d : std_logic := '0';
	
	signal bitvectord3196d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3196d : std_logic := '0';
	signal matchd3196d : std_logic := '0';
	
	signal bitvectord3197d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3197d : std_logic := '0';
	signal matchd3197d : std_logic := '0';
	
	signal bitvectord3198d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3198d : std_logic := '0';
	signal matchd3198d : std_logic := '0';
	
	signal bitvectord3199d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3199d : std_logic := '0';
	signal matchd3199d : std_logic := '0';
	
	signal bitvectord3200d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3200d : std_logic := '0';
	signal matchd3200d : std_logic := '0';
	
	signal bitvectord3201d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3201d : std_logic := '0';
	signal matchd3201d : std_logic := '0';
	
	signal bitvectord3202d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3202d : std_logic := '1';
	signal matchd3202d : std_logic := '0';
	
	signal bitvectord3203d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3203d : std_logic := '0';
	signal matchd3203d : std_logic := '0';
	
	signal bitvectord3204d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3204d : std_logic := '0';
	signal matchd3204d : std_logic := '0';
	
	signal bitvectord3205d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3205d : std_logic := '0';
	signal matchd3205d : std_logic := '0';
	
	signal bitvectord3206d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3206d : std_logic := '0';
	signal matchd3206d : std_logic := '0';
	
	signal bitvectord3207d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3207d : std_logic := '0';
	signal matchd3207d : std_logic := '0';
	
	signal bitvectord3208d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3208d : std_logic := '0';
	signal matchd3208d : std_logic := '0';
	
	signal bitvectord3209d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3209d : std_logic := '0';
	signal matchd3209d : std_logic := '0';
	
	signal bitvectord3210d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3210d : std_logic := '0';
	signal matchd3210d : std_logic := '0';
	
	signal bitvectord3211d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3211d : std_logic := '0';
	signal matchd3211d : std_logic := '0';
	
	signal bitvectord3212d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3212d : std_logic := '0';
	signal matchd3212d : std_logic := '0';
	
	signal bitvectord3213d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3213d : std_logic := '0';
	signal matchd3213d : std_logic := '0';
	
	signal bitvectord3214d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3214d : std_logic := '1';
	signal matchd3214d : std_logic := '0';
	
	signal bitvectord3215d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3215d : std_logic := '0';
	signal matchd3215d : std_logic := '0';
	
	signal bitvectord3216d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3216d : std_logic := '0';
	signal matchd3216d : std_logic := '0';
	
	signal bitvectord3217d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3217d : std_logic := '0';
	signal matchd3217d : std_logic := '0';
	
	signal bitvectord3218d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3218d : std_logic := '0';
	signal matchd3218d : std_logic := '0';
	
	signal bitvectord3219d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3219d : std_logic := '0';
	signal matchd3219d : std_logic := '0';
	
	signal bitvectord3220d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3220d : std_logic := '0';
	signal matchd3220d : std_logic := '0';
	
	signal bitvectord3221d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3221d : std_logic := '0';
	signal matchd3221d : std_logic := '0';
	
	signal bitvectord3222d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3222d : std_logic := '0';
	signal matchd3222d : std_logic := '0';
	
	signal bitvectord3223d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3223d : std_logic := '0';
	signal matchd3223d : std_logic := '0';
	
	signal bitvectord3224d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3224d : std_logic := '0';
	signal matchd3224d : std_logic := '0';
	
	signal bitvectord3225d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3225d : std_logic := '0';
	signal matchd3225d : std_logic := '0';
	
	signal bitvectord3226d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3226d : std_logic := '0';
	signal matchd3226d : std_logic := '0';
	
	signal bitvectord3227d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3227d : std_logic := '1';
	signal matchd3227d : std_logic := '0';
	
	signal bitvectord3228d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3228d : std_logic := '0';
	signal matchd3228d : std_logic := '0';
	
	signal bitvectord3229d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3229d : std_logic := '0';
	signal matchd3229d : std_logic := '0';
	
	signal bitvectord3230d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3230d : std_logic := '0';
	signal matchd3230d : std_logic := '0';
	
	signal bitvectord3231d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3231d : std_logic := '0';
	signal matchd3231d : std_logic := '0';
	
	signal bitvectord3232d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3232d : std_logic := '0';
	signal matchd3232d : std_logic := '0';
	
	signal bitvectord3233d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3233d : std_logic := '0';
	signal matchd3233d : std_logic := '0';
	
	signal bitvectord3234d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3234d : std_logic := '0';
	signal matchd3234d : std_logic := '0';
	
	signal bitvectord3235d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3235d : std_logic := '0';
	signal matchd3235d : std_logic := '0';
	
	signal bitvectord3236d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3236d : std_logic := '0';
	signal matchd3236d : std_logic := '0';
	
	signal bitvectord3237d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3237d : std_logic := '0';
	signal matchd3237d : std_logic := '0';
	
	signal bitvectord3238d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3238d : std_logic := '1';
	signal matchd3238d : std_logic := '0';
	
	signal bitvectord3239d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3239d : std_logic := '0';
	signal matchd3239d : std_logic := '0';
	
	signal bitvectord3240d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3240d : std_logic := '0';
	signal matchd3240d : std_logic := '0';
	
	signal bitvectord3241d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3241d : std_logic := '0';
	signal matchd3241d : std_logic := '0';
	
	signal bitvectord3242d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3242d : std_logic := '0';
	signal matchd3242d : std_logic := '0';
	
	signal bitvectord3243d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3243d : std_logic := '0';
	signal matchd3243d : std_logic := '0';
	
	signal bitvectord3244d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3244d : std_logic := '0';
	signal matchd3244d : std_logic := '0';
	
	signal bitvectord3245d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3245d : std_logic := '1';
	signal matchd3245d : std_logic := '0';
	
	signal bitvectord3246d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3246d : std_logic := '0';
	signal matchd3246d : std_logic := '0';
	
	signal bitvectord3247d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3247d : std_logic := '0';
	signal matchd3247d : std_logic := '0';
	
	signal bitvectord3248d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3248d : std_logic := '0';
	signal matchd3248d : std_logic := '0';
	
	signal bitvectord3249d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3249d : std_logic := '0';
	signal matchd3249d : std_logic := '0';
	
	signal bitvectord3250d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3250d : std_logic := '0';
	signal matchd3250d : std_logic := '0';
	
	signal bitvectord3251d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3251d : std_logic := '0';
	signal matchd3251d : std_logic := '0';
	
	signal bitvectord3252d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3252d : std_logic := '0';
	signal matchd3252d : std_logic := '0';
	
	signal bitvectord3253d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3253d : std_logic := '0';
	signal matchd3253d : std_logic := '0';
	
	signal bitvectord3254d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3254d : std_logic := '0';
	signal matchd3254d : std_logic := '0';
	
	signal bitvectord3255d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3255d : std_logic := '0';
	signal matchd3255d : std_logic := '0';
	
	signal bitvectord3256d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3256d : std_logic := '0';
	signal matchd3256d : std_logic := '0';
	
	signal bitvectord3257d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3257d : std_logic := '0';
	signal matchd3257d : std_logic := '0';
	
	signal bitvectord3258d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3258d : std_logic := '0';
	signal matchd3258d : std_logic := '0';
	
	signal bitvectord3259d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000";
	signal Enabled3259d : std_logic := '0';
	signal matchd3259d : std_logic := '0';
	
	signal bitvectord3260d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3260d : std_logic := '0';
	signal matchd3260d : std_logic := '0';
	
	signal bitvectord3261d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3261d : std_logic := '1';
	signal matchd3261d : std_logic := '0';
	
	signal bitvectord3262d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3262d : std_logic := '0';
	signal matchd3262d : std_logic := '0';
	
	signal bitvectord3263d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3263d : std_logic := '0';
	signal matchd3263d : std_logic := '0';
	
	signal bitvectord3264d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3264d : std_logic := '0';
	signal matchd3264d : std_logic := '0';
	
	signal bitvectord3265d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3265d : std_logic := '0';
	signal matchd3265d : std_logic := '0';
	
	signal bitvectord3266d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3266d : std_logic := '0';
	signal matchd3266d : std_logic := '0';
	
	signal bitvectord3267d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000";
	signal Enabled3267d : std_logic := '0';
	signal matchd3267d : std_logic := '0';
	
	signal bitvectord3268d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3268d : std_logic := '0';
	signal matchd3268d : std_logic := '0';
	
	signal bitvectord3269d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3269d : std_logic := '0';
	signal matchd3269d : std_logic := '0';
	
	signal bitvectord3270d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3270d : std_logic := '0';
	signal matchd3270d : std_logic := '0';
	
	signal bitvectord3271d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3271d : std_logic := '0';
	signal matchd3271d : std_logic := '0';
	
	signal bitvectord3272d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3272d : std_logic := '0';
	signal matchd3272d : std_logic := '0';
	
	signal bitvectord3273d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3273d : std_logic := '0';
	signal matchd3273d : std_logic := '0';
	
	signal bitvectord3274d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3274d : std_logic := '0';
	signal matchd3274d : std_logic := '0';
	
	signal bitvectord3275d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3275d : std_logic := '0';
	signal matchd3275d : std_logic := '0';
	
	signal bitvectord3276d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3276d : std_logic := '0';
	signal matchd3276d : std_logic := '0';
	
	signal bitvectord3277d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3277d : std_logic := '0';
	signal matchd3277d : std_logic := '0';
	
	signal bitvectord3278d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3278d : std_logic := '1';
	signal matchd3278d : std_logic := '0';
	
	signal bitvectord3279d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3279d : std_logic := '0';
	signal matchd3279d : std_logic := '0';
	
	signal bitvectord3280d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000";
	signal Enabled3280d : std_logic := '0';
	signal matchd3280d : std_logic := '0';
	
	signal bitvectord3281d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3281d : std_logic := '0';
	signal matchd3281d : std_logic := '0';
	
	signal bitvectord3282d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3282d : std_logic := '0';
	signal matchd3282d : std_logic := '0';
	
	signal bitvectord3283d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3283d : std_logic := '0';
	signal matchd3283d : std_logic := '0';
	
	signal bitvectord3284d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3284d : std_logic := '0';
	signal matchd3284d : std_logic := '0';
	
	signal bitvectord3285d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3285d : std_logic := '0';
	signal matchd3285d : std_logic := '0';
	
	signal bitvectord3286d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3286d : std_logic := '0';
	signal matchd3286d : std_logic := '0';
	
	signal bitvectord3287d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3287d : std_logic := '0';
	signal matchd3287d : std_logic := '0';
	
	signal bitvectord3288d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3288d : std_logic := '0';
	signal matchd3288d : std_logic := '0';
	
	signal bitvectord3289d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3289d : std_logic := '0';
	signal matchd3289d : std_logic := '0';
	
	signal bitvectord3290d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3290d : std_logic := '0';
	signal matchd3290d : std_logic := '0';
	
	signal bitvectord3291d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3291d : std_logic := '0';
	signal matchd3291d : std_logic := '0';
	
	signal bitvectord3292d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3292d : std_logic := '0';
	signal matchd3292d : std_logic := '0';
	
	signal bitvectord3293d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3293d : std_logic := '0';
	signal matchd3293d : std_logic := '0';
	
	signal bitvectord3294d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3294d : std_logic := '0';
	signal matchd3294d : std_logic := '0';
	
	signal bitvectord3296d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3296d : std_logic := '1';
	signal matchd3296d : std_logic := '0';
	
	signal bitvectord3297d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3297d : std_logic := '0';
	signal matchd3297d : std_logic := '0';
	
	signal bitvectord3298d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3298d : std_logic := '0';
	signal matchd3298d : std_logic := '0';
	
	signal bitvectord3299d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3299d : std_logic := '0';
	signal matchd3299d : std_logic := '0';
	
	signal bitvectord3300d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3300d : std_logic := '0';
	signal matchd3300d : std_logic := '0';
	
	signal bitvectord3301d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3301d : std_logic := '0';
	signal matchd3301d : std_logic := '0';
	
	signal bitvectord3302d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
	signal Enabled3302d : std_logic := '0';
	signal matchd3302d : std_logic := '0';
	
	signal bitvectord3303d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3303d : std_logic := '0';
	signal matchd3303d : std_logic := '0';
	
	signal bitvectord3304d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3304d : std_logic := '0';
	signal matchd3304d : std_logic := '0';
	
	signal bitvectord3305d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3305d : std_logic := '0';
	signal matchd3305d : std_logic := '0';
	
	signal bitvectord3306d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3306d : std_logic := '0';
	signal matchd3306d : std_logic := '0';
	
	signal bitvectord3307d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3307d : std_logic := '0';
	signal matchd3307d : std_logic := '0';
	
	signal bitvectord3308d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3308d : std_logic := '0';
	signal matchd3308d : std_logic := '0';
	
	signal bitvectord3309d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3309d : std_logic := '0';
	signal matchd3309d : std_logic := '0';
	
	signal bitvectord3310d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3310d : std_logic := '1';
	signal matchd3310d : std_logic := '0';
	
	signal bitvectord3311d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3311d : std_logic := '0';
	signal matchd3311d : std_logic := '0';
	
	signal bitvectord3312d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3312d : std_logic := '0';
	signal matchd3312d : std_logic := '0';
	
	signal bitvectord3313d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3313d : std_logic := '0';
	signal matchd3313d : std_logic := '0';
	
	signal bitvectord3314d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3314d : std_logic := '0';
	signal matchd3314d : std_logic := '0';
	
	signal bitvectord3315d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3315d : std_logic := '0';
	signal matchd3315d : std_logic := '0';
	
	signal bitvectord3316d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3316d : std_logic := '0';
	signal matchd3316d : std_logic := '0';
	
	signal bitvectord3317d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3317d : std_logic := '0';
	signal matchd3317d : std_logic := '0';
	
	signal bitvectord3318d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3318d : std_logic := '0';
	signal matchd3318d : std_logic := '0';
	
	signal bitvectord3319d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3319d : std_logic := '0';
	signal matchd3319d : std_logic := '0';
	
	signal bitvectord3320d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3320d : std_logic := '0';
	signal matchd3320d : std_logic := '0';
	
	signal bitvectord3321d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3321d : std_logic := '0';
	signal matchd3321d : std_logic := '0';
	
	signal bitvectord3322d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3322d : std_logic := '0';
	signal matchd3322d : std_logic := '0';
	
	signal bitvectord3323d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3323d : std_logic := '0';
	signal matchd3323d : std_logic := '0';
	
	signal bitvectord3324d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3324d : std_logic := '1';
	signal matchd3324d : std_logic := '0';
	
	signal bitvectord3325d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3325d : std_logic := '0';
	signal matchd3325d : std_logic := '0';
	
	signal bitvectord3326d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3326d : std_logic := '0';
	signal matchd3326d : std_logic := '0';
	
	signal bitvectord3327d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3327d : std_logic := '0';
	signal matchd3327d : std_logic := '0';
	
	signal bitvectord3328d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3328d : std_logic := '0';
	signal matchd3328d : std_logic := '0';
	
	signal bitvectord3329d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3329d : std_logic := '0';
	signal matchd3329d : std_logic := '0';
	
	signal bitvectord3330d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3330d : std_logic := '0';
	signal matchd3330d : std_logic := '0';
	
	signal bitvectord3331d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3331d : std_logic := '0';
	signal matchd3331d : std_logic := '0';
	
	signal bitvectord3332d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3332d : std_logic := '0';
	signal matchd3332d : std_logic := '0';
	
	signal bitvectord3333d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3333d : std_logic := '0';
	signal matchd3333d : std_logic := '0';
	
	signal bitvectord3334d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3334d : std_logic := '0';
	signal matchd3334d : std_logic := '0';
	
	signal bitvectord3335d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3335d : std_logic := '1';
	signal matchd3335d : std_logic := '0';
	
	signal bitvectord3336d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3336d : std_logic := '0';
	signal matchd3336d : std_logic := '0';
	
	signal bitvectord3337d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3337d : std_logic := '0';
	signal matchd3337d : std_logic := '0';
	
	signal bitvectord3338d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3338d : std_logic := '0';
	signal matchd3338d : std_logic := '0';
	
	signal bitvectord3339d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3339d : std_logic := '0';
	signal matchd3339d : std_logic := '0';
	
	signal bitvectord3340d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3340d : std_logic := '0';
	signal matchd3340d : std_logic := '0';
	
	signal bitvectord3341d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3341d : std_logic := '0';
	signal matchd3341d : std_logic := '0';
	
	signal bitvectord3342d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3342d : std_logic := '0';
	signal matchd3342d : std_logic := '0';
	
	signal bitvectord3343d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3343d : std_logic := '0';
	signal matchd3343d : std_logic := '0';
	
	signal bitvectord3344d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3344d : std_logic := '0';
	signal matchd3344d : std_logic := '0';
	
	signal bitvectord3345d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3345d : std_logic := '0';
	signal matchd3345d : std_logic := '0';
	
	signal bitvectord3346d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3346d : std_logic := '0';
	signal matchd3346d : std_logic := '0';
	
	signal bitvectord3347d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3347d : std_logic := '0';
	signal matchd3347d : std_logic := '0';
	
	signal bitvectord3348d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3348d : std_logic := '1';
	signal matchd3348d : std_logic := '0';
	
	signal bitvectord3349d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3349d : std_logic := '0';
	signal matchd3349d : std_logic := '0';
	
	signal bitvectord3350d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3350d : std_logic := '0';
	signal matchd3350d : std_logic := '0';
	
	signal bitvectord3351d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3351d : std_logic := '0';
	signal matchd3351d : std_logic := '0';
	
	signal bitvectord3352d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3352d : std_logic := '0';
	signal matchd3352d : std_logic := '0';
	
	signal bitvectord3353d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3353d : std_logic := '0';
	signal matchd3353d : std_logic := '0';
	
	signal bitvectord3354d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3354d : std_logic := '0';
	signal matchd3354d : std_logic := '0';
	
	signal bitvectord3355d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3355d : std_logic := '0';
	signal matchd3355d : std_logic := '0';
	
	signal bitvectord3356d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3356d : std_logic := '0';
	signal matchd3356d : std_logic := '0';
	
	signal bitvectord3357d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3357d : std_logic := '0';
	signal matchd3357d : std_logic := '0';
	
	signal bitvectord3358d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3358d : std_logic := '0';
	signal matchd3358d : std_logic := '0';
	
	signal bitvectord3359d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3359d : std_logic := '0';
	signal matchd3359d : std_logic := '0';
	
	signal bitvectord3360d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3360d : std_logic := '0';
	signal matchd3360d : std_logic := '0';
	
	signal bitvectord3361d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3361d : std_logic := '0';
	signal matchd3361d : std_logic := '0';
	
	signal bitvectord3362d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3362d : std_logic := '1';
	signal matchd3362d : std_logic := '0';
	
	signal bitvectord3363d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3363d : std_logic := '0';
	signal matchd3363d : std_logic := '0';
	
	signal bitvectord3364d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3364d : std_logic := '0';
	signal matchd3364d : std_logic := '0';
	
	signal bitvectord3365d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3365d : std_logic := '0';
	signal matchd3365d : std_logic := '0';
	
	signal bitvectord3366d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3366d : std_logic := '0';
	signal matchd3366d : std_logic := '0';
	
	signal bitvectord3367d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3367d : std_logic := '0';
	signal matchd3367d : std_logic := '0';
	
	signal bitvectord3368d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3368d : std_logic := '0';
	signal matchd3368d : std_logic := '0';
	
	signal bitvectord3369d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3369d : std_logic := '0';
	signal matchd3369d : std_logic := '0';
	
	signal bitvectord3370d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3370d : std_logic := '0';
	signal matchd3370d : std_logic := '0';
	
	signal bitvectord3371d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3371d : std_logic := '0';
	signal matchd3371d : std_logic := '0';
	
	signal bitvectord3372d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3372d : std_logic := '0';
	signal matchd3372d : std_logic := '0';
	
	signal bitvectord3373d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3373d : std_logic := '0';
	signal matchd3373d : std_logic := '0';
	
	signal bitvectord3374d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3374d : std_logic := '0';
	signal matchd3374d : std_logic := '0';
	
	signal bitvectord3375d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3375d : std_logic := '0';
	signal matchd3375d : std_logic := '0';
	
	signal bitvectord3376d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3376d : std_logic := '0';
	signal matchd3376d : std_logic := '0';
	
	signal bitvectord3377d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3377d : std_logic := '0';
	signal matchd3377d : std_logic := '0';
	
	signal bitvectord3378d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3378d : std_logic := '1';
	signal matchd3378d : std_logic := '0';
	
	signal bitvectord3379d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3379d : std_logic := '0';
	signal matchd3379d : std_logic := '0';
	
	signal bitvectord3380d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3380d : std_logic := '0';
	signal matchd3380d : std_logic := '0';
	
	signal bitvectord3381d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3381d : std_logic := '0';
	signal matchd3381d : std_logic := '0';
	
	signal bitvectord3382d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3382d : std_logic := '0';
	signal matchd3382d : std_logic := '0';
	
	signal bitvectord3383d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3383d : std_logic := '0';
	signal matchd3383d : std_logic := '0';
	
	signal bitvectord3384d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3384d : std_logic := '0';
	signal matchd3384d : std_logic := '0';
	
	signal bitvectord3385d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3385d : std_logic := '0';
	signal matchd3385d : std_logic := '0';
	
	signal bitvectord3386d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3386d : std_logic := '0';
	signal matchd3386d : std_logic := '0';
	
	signal bitvectord3387d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3387d : std_logic := '0';
	signal matchd3387d : std_logic := '0';
	
	signal bitvectord3388d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3388d : std_logic := '0';
	signal matchd3388d : std_logic := '0';
	
	signal bitvectord3389d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3389d : std_logic := '1';
	signal matchd3389d : std_logic := '0';
	
	signal bitvectord3390d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3390d : std_logic := '0';
	signal matchd3390d : std_logic := '0';
	
	signal bitvectord3391d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3391d : std_logic := '0';
	signal matchd3391d : std_logic := '0';
	
	signal bitvectord3392d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3392d : std_logic := '0';
	signal matchd3392d : std_logic := '0';
	
	signal bitvectord3393d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3393d : std_logic := '0';
	signal matchd3393d : std_logic := '0';
	
	signal bitvectord3394d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3394d : std_logic := '0';
	signal matchd3394d : std_logic := '0';
	
	signal bitvectord3395d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3395d : std_logic := '0';
	signal matchd3395d : std_logic := '0';
	
	signal bitvectord3396d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3396d : std_logic := '0';
	signal matchd3396d : std_logic := '0';
	
	signal bitvectord3397d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3397d : std_logic := '0';
	signal matchd3397d : std_logic := '0';
	
	signal bitvectord3398d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3398d : std_logic := '0';
	signal matchd3398d : std_logic := '0';
	
	signal bitvectord3399d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3399d : std_logic := '0';
	signal matchd3399d : std_logic := '0';
	
	signal bitvectord3400d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3400d : std_logic := '1';
	signal matchd3400d : std_logic := '0';
	
	signal bitvectord3401d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3401d : std_logic := '0';
	signal matchd3401d : std_logic := '0';
	
	signal bitvectord3402d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3402d : std_logic := '0';
	signal matchd3402d : std_logic := '0';
	
	signal bitvectord3403d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3403d : std_logic := '0';
	signal matchd3403d : std_logic := '0';
	
	signal bitvectord3404d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3404d : std_logic := '0';
	signal matchd3404d : std_logic := '0';
	
	signal bitvectord3405d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3405d : std_logic := '0';
	signal matchd3405d : std_logic := '0';
	
	signal bitvectord3406d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3406d : std_logic := '0';
	signal matchd3406d : std_logic := '0';
	
	signal bitvectord3407d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3407d : std_logic := '0';
	signal matchd3407d : std_logic := '0';
	
	signal bitvectord3408d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3408d : std_logic := '0';
	signal matchd3408d : std_logic := '0';
	
	signal bitvectord3409d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3409d : std_logic := '0';
	signal matchd3409d : std_logic := '0';
	
	signal bitvectord3410d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3410d : std_logic := '0';
	signal matchd3410d : std_logic := '0';
	
	signal bitvectord3411d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3411d : std_logic := '0';
	signal matchd3411d : std_logic := '0';
	
	signal bitvectord3412d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3412d : std_logic := '1';
	signal matchd3412d : std_logic := '0';
	
	signal bitvectord3413d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3413d : std_logic := '0';
	signal matchd3413d : std_logic := '0';
	
	signal bitvectord3414d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3414d : std_logic := '0';
	signal matchd3414d : std_logic := '0';
	
	signal bitvectord3415d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3415d : std_logic := '0';
	signal matchd3415d : std_logic := '0';
	
	signal bitvectord3416d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3416d : std_logic := '0';
	signal matchd3416d : std_logic := '0';
	
	signal bitvectord3417d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3417d : std_logic := '0';
	signal matchd3417d : std_logic := '0';
	
	signal bitvectord3418d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3418d : std_logic := '0';
	signal matchd3418d : std_logic := '0';
	
	signal bitvectord3419d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3419d : std_logic := '0';
	signal matchd3419d : std_logic := '0';
	
	signal bitvectord3420d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3420d : std_logic := '0';
	signal matchd3420d : std_logic := '0';
	
	signal bitvectord3421d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3421d : std_logic := '0';
	signal matchd3421d : std_logic := '0';
	
	signal bitvectord3422d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3422d : std_logic := '0';
	signal matchd3422d : std_logic := '0';
	
	signal bitvectord3423d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3423d : std_logic := '0';
	signal matchd3423d : std_logic := '0';
	
	signal bitvectord3424d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3424d : std_logic := '1';
	signal matchd3424d : std_logic := '0';
	
	signal bitvectord3425d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3425d : std_logic := '0';
	signal matchd3425d : std_logic := '0';
	
	signal bitvectord3426d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3426d : std_logic := '0';
	signal matchd3426d : std_logic := '0';
	
	signal bitvectord3427d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3427d : std_logic := '0';
	signal matchd3427d : std_logic := '0';
	
	signal bitvectord3428d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3428d : std_logic := '0';
	signal matchd3428d : std_logic := '0';
	
	signal bitvectord3429d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3429d : std_logic := '0';
	signal matchd3429d : std_logic := '0';
	
	signal bitvectord3430d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3430d : std_logic := '0';
	signal matchd3430d : std_logic := '0';
	
	signal bitvectord3431d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3431d : std_logic := '0';
	signal matchd3431d : std_logic := '0';
	
	signal bitvectord3432d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3432d : std_logic := '0';
	signal matchd3432d : std_logic := '0';
	
	signal bitvectord3433d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3433d : std_logic := '0';
	signal matchd3433d : std_logic := '0';
	
	signal bitvectord3434d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3434d : std_logic := '0';
	signal matchd3434d : std_logic := '0';
	
	signal bitvectord3435d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3435d : std_logic := '0';
	signal matchd3435d : std_logic := '0';
	
	signal bitvectord3436d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3436d : std_logic := '1';
	signal matchd3436d : std_logic := '0';
	
	signal bitvectord3437d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3437d : std_logic := '0';
	signal matchd3437d : std_logic := '0';
	
	signal bitvectord3438d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3438d : std_logic := '0';
	signal matchd3438d : std_logic := '0';
	
	signal bitvectord3439d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3439d : std_logic := '0';
	signal matchd3439d : std_logic := '0';
	
	signal bitvectord3440d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3440d : std_logic := '0';
	signal matchd3440d : std_logic := '0';
	
	signal bitvectord3441d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3441d : std_logic := '0';
	signal matchd3441d : std_logic := '0';
	
	signal bitvectord3442d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3442d : std_logic := '0';
	signal matchd3442d : std_logic := '0';
	
	signal bitvectord3443d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3443d : std_logic := '0';
	signal matchd3443d : std_logic := '0';
	
	signal bitvectord3444d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3444d : std_logic := '0';
	signal matchd3444d : std_logic := '0';
	
	signal bitvectord3445d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3445d : std_logic := '0';
	signal matchd3445d : std_logic := '0';
	
	signal bitvectord3446d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3446d : std_logic := '0';
	signal matchd3446d : std_logic := '0';
	
	signal bitvectord3447d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3447d : std_logic := '1';
	signal matchd3447d : std_logic := '0';
	
	signal bitvectord3448d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3448d : std_logic := '0';
	signal matchd3448d : std_logic := '0';
	
	signal bitvectord3449d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3449d : std_logic := '0';
	signal matchd3449d : std_logic := '0';
	
	signal bitvectord3450d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3450d : std_logic := '0';
	signal matchd3450d : std_logic := '0';
	
	signal bitvectord3451d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3451d : std_logic := '0';
	signal matchd3451d : std_logic := '0';
	
	signal bitvectord3452d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3452d : std_logic := '0';
	signal matchd3452d : std_logic := '0';
	
	signal bitvectord3453d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3453d : std_logic := '0';
	signal matchd3453d : std_logic := '0';
	
	signal bitvectord3454d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3454d : std_logic := '0';
	signal matchd3454d : std_logic := '0';
	
	signal bitvectord3455d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3455d : std_logic := '0';
	signal matchd3455d : std_logic := '0';
	
	signal bitvectord3456d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3456d : std_logic := '0';
	signal matchd3456d : std_logic := '0';
	
	signal bitvectord3457d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3457d : std_logic := '0';
	signal matchd3457d : std_logic := '0';
	
	signal bitvectord3458d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3458d : std_logic := '1';
	signal matchd3458d : std_logic := '0';
	
	signal bitvectord3459d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3459d : std_logic := '0';
	signal matchd3459d : std_logic := '0';
	
	signal bitvectord3460d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3460d : std_logic := '0';
	signal matchd3460d : std_logic := '0';
	
	signal bitvectord3461d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3461d : std_logic := '0';
	signal matchd3461d : std_logic := '0';
	
	signal bitvectord3462d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3462d : std_logic := '0';
	signal matchd3462d : std_logic := '0';
	
	signal bitvectord3463d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3463d : std_logic := '0';
	signal matchd3463d : std_logic := '0';
	
	signal bitvectord3464d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3464d : std_logic := '0';
	signal matchd3464d : std_logic := '0';
	
	signal bitvectord3465d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3465d : std_logic := '0';
	signal matchd3465d : std_logic := '0';
	
	signal bitvectord3466d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3466d : std_logic := '0';
	signal matchd3466d : std_logic := '0';
	
	signal bitvectord3467d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3467d : std_logic := '0';
	signal matchd3467d : std_logic := '0';
	
	signal bitvectord3468d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3468d : std_logic := '0';
	signal matchd3468d : std_logic := '0';
	
	signal bitvectord3469d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3469d : std_logic := '0';
	signal matchd3469d : std_logic := '0';
	
	signal bitvectord3470d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3470d : std_logic := '1';
	signal matchd3470d : std_logic := '0';
	
	signal bitvectord3471d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3471d : std_logic := '0';
	signal matchd3471d : std_logic := '0';
	
	signal bitvectord3472d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3472d : std_logic := '0';
	signal matchd3472d : std_logic := '0';
	
	signal bitvectord3473d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3473d : std_logic := '0';
	signal matchd3473d : std_logic := '0';
	
	signal bitvectord3474d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3474d : std_logic := '0';
	signal matchd3474d : std_logic := '0';
	
	signal bitvectord3475d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3475d : std_logic := '0';
	signal matchd3475d : std_logic := '0';
	
	signal bitvectord3476d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3476d : std_logic := '0';
	signal matchd3476d : std_logic := '0';
	
	signal bitvectord3477d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3477d : std_logic := '0';
	signal matchd3477d : std_logic := '0';
	
	signal bitvectord3478d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3478d : std_logic := '0';
	signal matchd3478d : std_logic := '0';
	
	signal bitvectord3479d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3479d : std_logic := '0';
	signal matchd3479d : std_logic := '0';
	
	signal bitvectord3480d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3480d : std_logic := '0';
	signal matchd3480d : std_logic := '0';
	
	signal bitvectord3481d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3481d : std_logic := '0';
	signal matchd3481d : std_logic := '0';
	
	signal bitvectord3482d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3482d : std_logic := '0';
	signal matchd3482d : std_logic := '0';
	
	signal bitvectord3483d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3483d : std_logic := '0';
	signal matchd3483d : std_logic := '0';
	
	signal bitvectord3484d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3484d : std_logic := '0';
	signal matchd3484d : std_logic := '0';
	
	signal bitvectord3485d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3485d : std_logic := '0';
	signal matchd3485d : std_logic := '0';
	
	signal bitvectord3486d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3486d : std_logic := '1';
	signal matchd3486d : std_logic := '0';
	
	signal bitvectord3487d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3487d : std_logic := '0';
	signal matchd3487d : std_logic := '0';
	
	signal bitvectord3488d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3488d : std_logic := '0';
	signal matchd3488d : std_logic := '0';
	
	signal bitvectord3489d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3489d : std_logic := '0';
	signal matchd3489d : std_logic := '0';
	
	signal bitvectord3490d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3490d : std_logic := '0';
	signal matchd3490d : std_logic := '0';
	
	signal bitvectord3491d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3491d : std_logic := '0';
	signal matchd3491d : std_logic := '0';
	
	signal bitvectord3492d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3492d : std_logic := '0';
	signal matchd3492d : std_logic := '0';
	
	signal bitvectord3493d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3493d : std_logic := '0';
	signal matchd3493d : std_logic := '0';
	
	signal bitvectord3494d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3494d : std_logic := '0';
	signal matchd3494d : std_logic := '0';
	
	signal bitvectord3495d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3495d : std_logic := '0';
	signal matchd3495d : std_logic := '0';
	
	signal bitvectord3496d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3496d : std_logic := '0';
	signal matchd3496d : std_logic := '0';
	
	signal bitvectord3497d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3497d : std_logic := '0';
	signal matchd3497d : std_logic := '0';
	
	signal bitvectord3498d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3498d : std_logic := '0';
	signal matchd3498d : std_logic := '0';
	
	signal bitvectord3499d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3499d : std_logic := '0';
	signal matchd3499d : std_logic := '0';
	
	signal bitvectord3500d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3500d : std_logic := '0';
	signal matchd3500d : std_logic := '0';
	
	signal bitvectord3501d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3501d : std_logic := '0';
	signal matchd3501d : std_logic := '0';
	
	signal bitvectord3502d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3502d : std_logic := '0';
	signal matchd3502d : std_logic := '0';
	
	signal bitvectord3503d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3503d : std_logic := '1';
	signal matchd3503d : std_logic := '0';
	
	signal bitvectord3504d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3504d : std_logic := '0';
	signal matchd3504d : std_logic := '0';
	
	signal bitvectord3505d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3505d : std_logic := '0';
	signal matchd3505d : std_logic := '0';
	
	signal bitvectord3506d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3506d : std_logic := '0';
	signal matchd3506d : std_logic := '0';
	
	signal bitvectord3507d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3507d : std_logic := '0';
	signal matchd3507d : std_logic := '0';
	
	signal bitvectord3508d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3508d : std_logic := '0';
	signal matchd3508d : std_logic := '0';
	
	signal bitvectord3509d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3509d : std_logic := '0';
	signal matchd3509d : std_logic := '0';
	
	signal bitvectord3510d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3510d : std_logic := '0';
	signal matchd3510d : std_logic := '0';
	
	signal bitvectord3511d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3511d : std_logic := '0';
	signal matchd3511d : std_logic := '0';
	
	signal bitvectord3512d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3512d : std_logic := '0';
	signal matchd3512d : std_logic := '0';
	
	signal bitvectord3513d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3513d : std_logic := '0';
	signal matchd3513d : std_logic := '0';
	
	signal bitvectord3514d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3514d : std_logic := '0';
	signal matchd3514d : std_logic := '0';
	
	signal bitvectord3515d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3515d : std_logic := '0';
	signal matchd3515d : std_logic := '0';
	
	signal bitvectord3516d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3516d : std_logic := '0';
	signal matchd3516d : std_logic := '0';
	
	signal bitvectord3517d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3517d : std_logic := '0';
	signal matchd3517d : std_logic := '0';
	
	signal bitvectord3518d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3518d : std_logic := '0';
	signal matchd3518d : std_logic := '0';
	
	signal bitvectord3519d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3519d : std_logic := '0';
	signal matchd3519d : std_logic := '0';
	
	signal bitvectord3520d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3520d : std_logic := '1';
	signal matchd3520d : std_logic := '0';
	
	signal bitvectord3521d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3521d : std_logic := '0';
	signal matchd3521d : std_logic := '0';
	
	signal bitvectord3522d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3522d : std_logic := '0';
	signal matchd3522d : std_logic := '0';
	
	signal bitvectord3523d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3523d : std_logic := '0';
	signal matchd3523d : std_logic := '0';
	
	signal bitvectord3524d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3524d : std_logic := '0';
	signal matchd3524d : std_logic := '0';
	
	signal bitvectord3525d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3525d : std_logic := '0';
	signal matchd3525d : std_logic := '0';
	
	signal bitvectord3526d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3526d : std_logic := '0';
	signal matchd3526d : std_logic := '0';
	
	signal bitvectord3527d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3527d : std_logic := '0';
	signal matchd3527d : std_logic := '0';
	
	signal bitvectord3528d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3528d : std_logic := '0';
	signal matchd3528d : std_logic := '0';
	
	signal bitvectord3529d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3529d : std_logic := '0';
	signal matchd3529d : std_logic := '0';
	
	signal bitvectord3530d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3530d : std_logic := '0';
	signal matchd3530d : std_logic := '0';
	
	signal bitvectord3531d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3531d : std_logic := '0';
	signal matchd3531d : std_logic := '0';
	
	signal bitvectord3532d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3532d : std_logic := '0';
	signal matchd3532d : std_logic := '0';
	
	signal bitvectord3533d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3533d : std_logic := '0';
	signal matchd3533d : std_logic := '0';
	
	signal bitvectord3534d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3534d : std_logic := '0';
	signal matchd3534d : std_logic := '0';
	
	signal bitvectord3535d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3535d : std_logic := '0';
	signal matchd3535d : std_logic := '0';
	
	signal bitvectord3536d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3536d : std_logic := '0';
	signal matchd3536d : std_logic := '0';
	
	signal bitvectord3537d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3537d : std_logic := '0';
	signal matchd3537d : std_logic := '0';
	
	signal bitvectord3538d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3538d : std_logic := '0';
	signal matchd3538d : std_logic := '0';
	
	signal bitvectord3539d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3539d : std_logic := '0';
	signal matchd3539d : std_logic := '0';
	
	signal bitvectord3540d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3540d : std_logic := '0';
	signal matchd3540d : std_logic := '0';
	
	signal bitvectord3541d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3541d : std_logic := '0';
	signal matchd3541d : std_logic := '0';
	
	signal bitvectord3542d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3542d : std_logic := '1';
	signal matchd3542d : std_logic := '0';
	
	signal bitvectord3543d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3543d : std_logic := '0';
	signal matchd3543d : std_logic := '0';
	
	signal bitvectord3544d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3544d : std_logic := '0';
	signal matchd3544d : std_logic := '0';
	
	signal bitvectord3545d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3545d : std_logic := '0';
	signal matchd3545d : std_logic := '0';
	
	signal bitvectord3546d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3546d : std_logic := '0';
	signal matchd3546d : std_logic := '0';
	
	signal bitvectord3547d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3547d : std_logic := '0';
	signal matchd3547d : std_logic := '0';
	
	signal bitvectord3548d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3548d : std_logic := '0';
	signal matchd3548d : std_logic := '0';
	
	signal bitvectord3549d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3549d : std_logic := '0';
	signal matchd3549d : std_logic := '0';
	
	signal bitvectord3550d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3550d : std_logic := '0';
	signal matchd3550d : std_logic := '0';
	
	signal bitvectord3551d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3551d : std_logic := '0';
	signal matchd3551d : std_logic := '0';
	
	signal bitvectord3552d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3552d : std_logic := '0';
	signal matchd3552d : std_logic := '0';
	
	signal bitvectord3553d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3553d : std_logic := '0';
	signal matchd3553d : std_logic := '0';
	
	signal bitvectord3554d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3554d : std_logic := '0';
	signal matchd3554d : std_logic := '0';
	
	signal bitvectord3555d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3555d : std_logic := '0';
	signal matchd3555d : std_logic := '0';
	
	signal bitvectord3556d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3556d : std_logic := '0';
	signal matchd3556d : std_logic := '0';
	
	signal bitvectord3557d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3557d : std_logic := '0';
	signal matchd3557d : std_logic := '0';
	
	signal bitvectord3558d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3558d : std_logic := '1';
	signal matchd3558d : std_logic := '0';
	
	signal bitvectord3559d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3559d : std_logic := '0';
	signal matchd3559d : std_logic := '0';
	
	signal bitvectord3560d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3560d : std_logic := '0';
	signal matchd3560d : std_logic := '0';
	
	signal bitvectord3561d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3561d : std_logic := '0';
	signal matchd3561d : std_logic := '0';
	
	signal bitvectord3562d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3562d : std_logic := '0';
	signal matchd3562d : std_logic := '0';
	
	signal bitvectord3563d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3563d : std_logic := '0';
	signal matchd3563d : std_logic := '0';
	
	signal bitvectord3564d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3564d : std_logic := '0';
	signal matchd3564d : std_logic := '0';
	
	signal bitvectord3565d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3565d : std_logic := '0';
	signal matchd3565d : std_logic := '0';
	
	signal bitvectord3566d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3566d : std_logic := '0';
	signal matchd3566d : std_logic := '0';
	
	signal bitvectord3567d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3567d : std_logic := '0';
	signal matchd3567d : std_logic := '0';
	
	signal bitvectord3568d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3568d : std_logic := '0';
	signal matchd3568d : std_logic := '0';
	
	signal bitvectord3569d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3569d : std_logic := '0';
	signal matchd3569d : std_logic := '0';
	
	signal bitvectord3570d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3570d : std_logic := '0';
	signal matchd3570d : std_logic := '0';
	
	signal bitvectord3571d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3571d : std_logic := '0';
	signal matchd3571d : std_logic := '0';
	
	signal bitvectord3572d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3572d : std_logic := '0';
	signal matchd3572d : std_logic := '0';
	
	signal bitvectord3573d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3573d : std_logic := '0';
	signal matchd3573d : std_logic := '0';
	
	signal bitvectord3574d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3574d : std_logic := '0';
	signal matchd3574d : std_logic := '0';
	
	signal bitvectord3575d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3575d : std_logic := '0';
	signal matchd3575d : std_logic := '0';
	
	signal bitvectord3576d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000";
	signal Enabled3576d : std_logic := '0';
	signal matchd3576d : std_logic := '0';
	
	signal bitvectord3577d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3577d : std_logic := '0';
	signal matchd3577d : std_logic := '0';
	
	signal bitvectord3578d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3578d : std_logic := '1';
	signal matchd3578d : std_logic := '0';
	
	signal bitvectord3579d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3579d : std_logic := '0';
	signal matchd3579d : std_logic := '0';
	
	signal bitvectord3580d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3580d : std_logic := '0';
	signal matchd3580d : std_logic := '0';
	
	signal bitvectord3581d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3581d : std_logic := '0';
	signal matchd3581d : std_logic := '0';
	
	signal bitvectord3582d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3582d : std_logic := '0';
	signal matchd3582d : std_logic := '0';
	
	signal bitvectord3583d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3583d : std_logic := '0';
	signal matchd3583d : std_logic := '0';
	
	signal bitvectord3584d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3584d : std_logic := '0';
	signal matchd3584d : std_logic := '0';
	
	signal bitvectord3585d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3585d : std_logic := '0';
	signal matchd3585d : std_logic := '0';
	
	signal bitvectord3586d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3586d : std_logic := '0';
	signal matchd3586d : std_logic := '0';
	
	signal bitvectord3587d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3587d : std_logic := '0';
	signal matchd3587d : std_logic := '0';
	
	signal bitvectord3588d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3588d : std_logic := '0';
	signal matchd3588d : std_logic := '0';
	
	signal bitvectord3589d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3589d : std_logic := '0';
	signal matchd3589d : std_logic := '0';
	
	signal bitvectord3590d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3590d : std_logic := '0';
	signal matchd3590d : std_logic := '0';
	
	signal bitvectord3591d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3591d : std_logic := '0';
	signal matchd3591d : std_logic := '0';
	
	signal bitvectord3592d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3592d : std_logic := '0';
	signal matchd3592d : std_logic := '0';
	
	signal bitvectord3593d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3593d : std_logic := '0';
	signal matchd3593d : std_logic := '0';
	
	signal bitvectord3594d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3594d : std_logic := '0';
	signal matchd3594d : std_logic := '0';
	
	signal bitvectord3595d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3595d : std_logic := '1';
	signal matchd3595d : std_logic := '0';
	
	signal bitvectord3596d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3596d : std_logic := '0';
	signal matchd3596d : std_logic := '0';
	
	signal bitvectord3597d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3597d : std_logic := '0';
	signal matchd3597d : std_logic := '0';
	
	signal bitvectord3598d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3598d : std_logic := '0';
	signal matchd3598d : std_logic := '0';
	
	signal bitvectord3599d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3599d : std_logic := '0';
	signal matchd3599d : std_logic := '0';
	
	signal bitvectord3600d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3600d : std_logic := '0';
	signal matchd3600d : std_logic := '0';
	
	signal bitvectord3601d : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111";
	signal Enabled3601d : std_logic := '0';
	signal matchd3601d : std_logic := '0';
	
	signal bitvectord3602d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
	signal Enabled3602d : std_logic := '0';
	signal matchd3602d : std_logic := '0';
	
	signal bitvectord3603d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3603d : std_logic := '0';
	signal matchd3603d : std_logic := '0';
	
	signal bitvectord3604d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enabled3604d : std_logic := '0';
	signal matchd3604d : std_logic := '0';
	
	signal bitvectord3605d : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
	signal Enabled3605d : std_logic := '0';
	signal matchd3605d : std_logic := '0';
	
	--- ORs
	signal matchd269d : std_logic := '0';
	
	signal matchd313d : std_logic := '0';
	
	signal matchd356d : std_logic := '0';
	
	signal matchd433d : std_logic := '0';
	
	signal matchd505d : std_logic := '0';
	
	signal matchd554d : std_logic := '0';
	
	signal matchd626d : std_logic := '0';
	
	signal matchd725d : std_logic := '0';
	
	signal matchd818d : std_logic := '0';
	
	signal matchd906d : std_logic := '0';
	
	signal matchd985d : std_logic := '0';
	
	signal matchd1119d : std_logic := '0';
	
	signal matchd1299d : std_logic := '0';
	
	signal matchd1763d : std_logic := '0';
	
	signal matchd1851d : std_logic := '0';
	
	signal matchd2324d : std_logic := '0';
	
	signal matchd2397d : std_logic := '0';
	
	signal matchd2836d : std_logic := '0';
	
	signal matchd2869d : std_logic := '0';
	
	signal matchd3058d : std_logic := '0';
	
	signal matchd3116d : std_logic := '0';
	
	signal matchd3182d : std_logic := '0';
	
	signal matchd3295d : std_logic := '0';
	
	
	--- ANDs
	
	--- Counters


begin
	--- STEs
	-- d2d
	sted2d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2d,
			Enable=>Enabled2d,
			match=>matchd2d,
			run=>run);

	-- d3d
	sted3d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3d,
			Enable=>Enabled3d,
			match=>matchd3d,
			run=>run);

	Enabled3d <= matchd2d;
	-- d4d
	sted4d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord4d,
			Enable=>Enabled4d,
			match=>matchd4d,
			run=>run);

	Enabled4d <= matchd3d;
	-- d5d
	sted5d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord5d,
			Enable=>Enabled5d,
			match=>matchd5d,
			run=>run);

	Enabled5d <= matchd4d;
	-- d6d
	sted6d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord6d,
			Enable=>Enabled6d,
			match=>matchd6d,
			run=>run);

	Enabled6d <= matchd5d;
	-- d7d
	sted7d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord7d,
			Enable=>Enabled7d,
			match=>matchd7d,
			run=>run);

	Enabled7d <= matchd6d;
	-- d8d
	sted8d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord8d,
			Enable=>Enabled8d,
			match=>matchd8d,
			run=>run);

	Enabled8d <= matchd7d;
	-- d9d
	sted9d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord9d,
			Enable=>Enabled9d,
			match=>matchd9d,
			run=>run);

	Enabled9d <= matchd8d;
	-- d10d
	sted10d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord10d,
			Enable=>Enabled10d,
			match=>matchd10d,
			run=>run);

	Enabled10d <= matchd9d;
	-- d11d
	sted11d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord11d,
			Enable=>Enabled11d,
			match=>matchd11d,
			run=>run);

	Enabled11d <= matchd10d;
	-- d12d
	sted12d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord12d,
			Enable=>Enabled12d,
			match=>matchd12d,
			run=>run);

	Enabled12d <= matchd11d;
	-- d13d
	sted13d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord13d,
			Enable=>Enabled13d,
			match=>matchd13d,
			run=>run);

	Enabled13d <= matchd12d;
	-- d14d
	sted14d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord14d,
			Enable=>Enabled14d,
			match=>matchd14d,
			run=>run);

	Enabled14d <= matchd13d;
	-- d15d
	sted15d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord15d,
			Enable=>Enabled15d,
			match=>matchd15d,
			run=>run);

	Enabled15d <= matchd15d OR matchd14d;
	-- d16d
	sted16d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord16d,
			Enable=>Enabled16d,
			match=>matchd16d,
			run=>run);

	reports(0) <= matchd16d;
	Enabled16d <= matchd15d;
	-- d17d
	sted17d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord17d,
			Enable=>Enabled17d,
			match=>matchd17d,
			run=>run);

	-- d18d
	sted18d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord18d,
			Enable=>Enabled18d,
			match=>matchd18d,
			run=>run);

	Enabled18d <= matchd17d;
	-- d19d
	sted19d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord19d,
			Enable=>Enabled19d,
			match=>matchd19d,
			run=>run);

	Enabled19d <= matchd18d;
	-- d20d
	sted20d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord20d,
			Enable=>Enabled20d,
			match=>matchd20d,
			run=>run);

	Enabled20d <= matchd19d;
	-- d21d
	sted21d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord21d,
			Enable=>Enabled21d,
			match=>matchd21d,
			run=>run);

	Enabled21d <= matchd20d;
	-- d22d
	sted22d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord22d,
			Enable=>Enabled22d,
			match=>matchd22d,
			run=>run);

	Enabled22d <= matchd21d OR matchd22d;
	-- d23d
	sted23d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord23d,
			Enable=>Enabled23d,
			match=>matchd23d,
			run=>run);

	Enabled23d <= matchd22d;
	-- d24d
	sted24d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord24d,
			Enable=>Enabled24d,
			match=>matchd24d,
			run=>run);

	Enabled24d <= matchd23d;
	-- d25d
	sted25d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord25d,
			Enable=>Enabled25d,
			match=>matchd25d,
			run=>run);

	Enabled25d <= matchd24d;
	-- d26d
	sted26d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord26d,
			Enable=>Enabled26d,
			match=>matchd26d,
			run=>run);

	Enabled26d <= matchd25d;
	-- d27d
	sted27d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord27d,
			Enable=>Enabled27d,
			match=>matchd27d,
			run=>run);

	Enabled27d <= matchd26d;
	-- d28d
	sted28d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord28d,
			Enable=>Enabled28d,
			match=>matchd28d,
			run=>run);

	Enabled28d <= matchd27d;
	-- d29d
	sted29d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord29d,
			Enable=>Enabled29d,
			match=>matchd29d,
			run=>run);

	Enabled29d <= matchd28d;
	-- d30d
	sted30d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord30d,
			Enable=>Enabled30d,
			match=>matchd30d,
			run=>run);

	Enabled30d <= matchd29d;
	-- d31d
	sted31d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord31d,
			Enable=>Enabled31d,
			match=>matchd31d,
			run=>run);

	reports(1) <= matchd31d;
	Enabled31d <= matchd30d;
	-- d32d
	sted32d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord32d,
			Enable=>Enabled32d,
			match=>matchd32d,
			run=>run);

	-- d33d
	sted33d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord33d,
			Enable=>Enabled33d,
			match=>matchd33d,
			run=>run);

	Enabled33d <= matchd32d OR matchd33d;
	-- d34d
	sted34d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord34d,
			Enable=>Enabled34d,
			match=>matchd34d,
			run=>run);

	Enabled34d <= matchd33d;
	-- d35d
	sted35d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord35d,
			Enable=>Enabled35d,
			match=>matchd35d,
			run=>run);

	Enabled35d <= matchd34d;
	-- d36d
	sted36d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord36d,
			Enable=>Enabled36d,
			match=>matchd36d,
			run=>run);

	Enabled36d <= matchd35d;
	-- d37d
	sted37d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord37d,
			Enable=>Enabled37d,
			match=>matchd37d,
			run=>run);

	Enabled37d <= matchd36d;
	-- d38d
	sted38d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord38d,
			Enable=>Enabled38d,
			match=>matchd38d,
			run=>run);

	Enabled38d <= matchd37d;
	-- d39d
	sted39d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord39d,
			Enable=>Enabled39d,
			match=>matchd39d,
			run=>run);

	Enabled39d <= matchd38d;
	-- d40d
	sted40d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord40d,
			Enable=>Enabled40d,
			match=>matchd40d,
			run=>run);

	Enabled40d <= matchd39d;
	-- d41d
	sted41d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord41d,
			Enable=>Enabled41d,
			match=>matchd41d,
			run=>run);

	Enabled41d <= matchd40d;
	-- d42d
	sted42d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord42d,
			Enable=>Enabled42d,
			match=>matchd42d,
			run=>run);

	Enabled42d <= matchd41d;
	-- d43d
	sted43d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord43d,
			Enable=>Enabled43d,
			match=>matchd43d,
			run=>run);

	Enabled43d <= matchd42d;
	-- d44d
	sted44d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord44d,
			Enable=>Enabled44d,
			match=>matchd44d,
			run=>run);

	Enabled44d <= matchd43d;
	-- d45d
	sted45d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord45d,
			Enable=>Enabled45d,
			match=>matchd45d,
			run=>run);

	Enabled45d <= matchd45d OR matchd44d;
	-- d46d
	sted46d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord46d,
			Enable=>Enabled46d,
			match=>matchd46d,
			run=>run);

	reports(2) <= matchd46d;
	Enabled46d <= matchd45d;
	-- d47d
	sted47d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord47d,
			Enable=>Enabled47d,
			match=>matchd47d,
			run=>run);

	-- d48d
	sted48d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord48d,
			Enable=>Enabled48d,
			match=>matchd48d,
			run=>run);

	Enabled48d <= matchd47d;
	-- d49d
	sted49d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord49d,
			Enable=>Enabled49d,
			match=>matchd49d,
			run=>run);

	Enabled49d <= matchd48d;
	-- d50d
	sted50d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord50d,
			Enable=>Enabled50d,
			match=>matchd50d,
			run=>run);

	Enabled50d <= matchd49d OR matchd50d;
	-- d51d
	sted51d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord51d,
			Enable=>Enabled51d,
			match=>matchd51d,
			run=>run);

	Enabled51d <= matchd50d;
	-- d52d
	sted52d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord52d,
			Enable=>Enabled52d,
			match=>matchd52d,
			run=>run);

	Enabled52d <= matchd51d;
	-- d53d
	sted53d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord53d,
			Enable=>Enabled53d,
			match=>matchd53d,
			run=>run);

	Enabled53d <= matchd52d;
	-- d54d
	sted54d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord54d,
			Enable=>Enabled54d,
			match=>matchd54d,
			run=>run);

	Enabled54d <= matchd53d;
	-- d55d
	sted55d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord55d,
			Enable=>Enabled55d,
			match=>matchd55d,
			run=>run);

	Enabled55d <= matchd54d;
	-- d56d
	sted56d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord56d,
			Enable=>Enabled56d,
			match=>matchd56d,
			run=>run);

	Enabled56d <= matchd55d;
	-- d57d
	sted57d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord57d,
			Enable=>Enabled57d,
			match=>matchd57d,
			run=>run);

	Enabled57d <= matchd56d;
	-- d58d
	sted58d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord58d,
			Enable=>Enabled58d,
			match=>matchd58d,
			run=>run);

	Enabled58d <= matchd57d;
	-- d59d
	sted59d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord59d,
			Enable=>Enabled59d,
			match=>matchd59d,
			run=>run);

	reports(3) <= matchd59d;
	Enabled59d <= matchd58d;
	-- d60d
	sted60d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord60d,
			Enable=>Enabled60d,
			match=>matchd60d,
			run=>run);

	-- d61d
	sted61d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord61d,
			Enable=>Enabled61d,
			match=>matchd61d,
			run=>run);

	Enabled61d <= matchd60d OR matchd61d;
	-- d62d
	sted62d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord62d,
			Enable=>Enabled62d,
			match=>matchd62d,
			run=>run);

	Enabled62d <= matchd61d;
	-- d63d
	sted63d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord63d,
			Enable=>Enabled63d,
			match=>matchd63d,
			run=>run);

	Enabled63d <= matchd62d;
	-- d64d
	sted64d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord64d,
			Enable=>Enabled64d,
			match=>matchd64d,
			run=>run);

	Enabled64d <= matchd63d;
	-- d65d
	sted65d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord65d,
			Enable=>Enabled65d,
			match=>matchd65d,
			run=>run);

	Enabled65d <= matchd64d;
	-- d66d
	sted66d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord66d,
			Enable=>Enabled66d,
			match=>matchd66d,
			run=>run);

	Enabled66d <= matchd65d;
	-- d67d
	sted67d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord67d,
			Enable=>Enabled67d,
			match=>matchd67d,
			run=>run);

	Enabled67d <= matchd66d;
	-- d68d
	sted68d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord68d,
			Enable=>Enabled68d,
			match=>matchd68d,
			run=>run);

	Enabled68d <= matchd67d;
	-- d69d
	sted69d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord69d,
			Enable=>Enabled69d,
			match=>matchd69d,
			run=>run);

	Enabled69d <= matchd68d;
	-- d70d
	sted70d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord70d,
			Enable=>Enabled70d,
			match=>matchd70d,
			run=>run);

	Enabled70d <= matchd69d OR matchd70d;
	-- d71d
	sted71d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord71d,
			Enable=>Enabled71d,
			match=>matchd71d,
			run=>run);

	reports(4) <= matchd71d;
	Enabled71d <= matchd70d;
	-- d72d
	sted72d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord72d,
			Enable=>Enabled72d,
			match=>matchd72d,
			run=>run);

	-- d73d
	sted73d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord73d,
			Enable=>Enabled73d,
			match=>matchd73d,
			run=>run);

	Enabled73d <= matchd72d;
	-- d74d
	sted74d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord74d,
			Enable=>Enabled74d,
			match=>matchd74d,
			run=>run);

	Enabled74d <= matchd73d;
	-- d75d
	sted75d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord75d,
			Enable=>Enabled75d,
			match=>matchd75d,
			run=>run);

	Enabled75d <= matchd74d;
	-- d76d
	sted76d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord76d,
			Enable=>Enabled76d,
			match=>matchd76d,
			run=>run);

	Enabled76d <= matchd75d;
	-- d77d
	sted77d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord77d,
			Enable=>Enabled77d,
			match=>matchd77d,
			run=>run);

	Enabled77d <= matchd76d;
	-- d78d
	sted78d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord78d,
			Enable=>Enabled78d,
			match=>matchd78d,
			run=>run);

	Enabled78d <= matchd77d;
	-- d79d
	sted79d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord79d,
			Enable=>Enabled79d,
			match=>matchd79d,
			run=>run);

	Enabled79d <= matchd78d;
	-- d80d
	sted80d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord80d,
			Enable=>Enabled80d,
			match=>matchd80d,
			run=>run);

	Enabled80d <= matchd79d;
	-- d81d
	sted81d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord81d,
			Enable=>Enabled81d,
			match=>matchd81d,
			run=>run);

	Enabled81d <= matchd80d;
	-- d82d
	sted82d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord82d,
			Enable=>Enabled82d,
			match=>matchd82d,
			run=>run);

	Enabled82d <= matchd81d;
	-- d83d
	sted83d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord83d,
			Enable=>Enabled83d,
			match=>matchd83d,
			run=>run);

	Enabled83d <= matchd82d;
	-- d84d
	sted84d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord84d,
			Enable=>Enabled84d,
			match=>matchd84d,
			run=>run);

	Enabled84d <= matchd83d OR matchd84d;
	-- d85d
	sted85d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord85d,
			Enable=>Enabled85d,
			match=>matchd85d,
			run=>run);

	reports(5) <= matchd85d;
	Enabled85d <= matchd84d;
	-- d86d
	sted86d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord86d,
			Enable=>Enabled86d,
			match=>matchd86d,
			run=>run);

	-- d87d
	sted87d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord87d,
			Enable=>Enabled87d,
			match=>matchd87d,
			run=>run);

	Enabled87d <= matchd86d OR matchd87d;
	-- d88d
	sted88d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord88d,
			Enable=>Enabled88d,
			match=>matchd88d,
			run=>run);

	Enabled88d <= matchd87d;
	-- d89d
	sted89d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord89d,
			Enable=>Enabled89d,
			match=>matchd89d,
			run=>run);

	Enabled89d <= matchd88d;
	-- d90d
	sted90d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord90d,
			Enable=>Enabled90d,
			match=>matchd90d,
			run=>run);

	Enabled90d <= matchd89d;
	-- d91d
	sted91d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord91d,
			Enable=>Enabled91d,
			match=>matchd91d,
			run=>run);

	Enabled91d <= matchd90d;
	-- d92d
	sted92d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord92d,
			Enable=>Enabled92d,
			match=>matchd92d,
			run=>run);

	Enabled92d <= matchd91d;
	-- d93d
	sted93d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord93d,
			Enable=>Enabled93d,
			match=>matchd93d,
			run=>run);

	Enabled93d <= matchd92d;
	-- d94d
	sted94d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord94d,
			Enable=>Enabled94d,
			match=>matchd94d,
			run=>run);

	Enabled94d <= matchd93d;
	-- d95d
	sted95d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord95d,
			Enable=>Enabled95d,
			match=>matchd95d,
			run=>run);

	Enabled95d <= matchd94d;
	-- d96d
	sted96d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord96d,
			Enable=>Enabled96d,
			match=>matchd96d,
			run=>run);

	Enabled96d <= matchd95d;
	-- d97d
	sted97d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord97d,
			Enable=>Enabled97d,
			match=>matchd97d,
			run=>run);

	Enabled97d <= matchd96d;
	-- d98d
	sted98d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord98d,
			Enable=>Enabled98d,
			match=>matchd98d,
			run=>run);

	Enabled98d <= matchd98d OR matchd97d;
	-- d99d
	sted99d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord99d,
			Enable=>Enabled99d,
			match=>matchd99d,
			run=>run);

	reports(6) <= matchd99d;
	Enabled99d <= matchd98d;
	-- d100d
	sted100d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord100d,
			Enable=>Enabled100d,
			match=>matchd100d,
			run=>run);

	-- d101d
	sted101d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord101d,
			Enable=>Enabled101d,
			match=>matchd101d,
			run=>run);

	Enabled101d <= matchd101d OR matchd100d;
	-- d102d
	sted102d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord102d,
			Enable=>Enabled102d,
			match=>matchd102d,
			run=>run);

	Enabled102d <= matchd101d;
	-- d103d
	sted103d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord103d,
			Enable=>Enabled103d,
			match=>matchd103d,
			run=>run);

	Enabled103d <= matchd102d;
	-- d104d
	sted104d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord104d,
			Enable=>Enabled104d,
			match=>matchd104d,
			run=>run);

	Enabled104d <= matchd103d;
	-- d105d
	sted105d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord105d,
			Enable=>Enabled105d,
			match=>matchd105d,
			run=>run);

	Enabled105d <= matchd104d;
	-- d106d
	sted106d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord106d,
			Enable=>Enabled106d,
			match=>matchd106d,
			run=>run);

	Enabled106d <= matchd105d;
	-- d107d
	sted107d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord107d,
			Enable=>Enabled107d,
			match=>matchd107d,
			run=>run);

	Enabled107d <= matchd106d;
	-- d108d
	sted108d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord108d,
			Enable=>Enabled108d,
			match=>matchd108d,
			run=>run);

	Enabled108d <= matchd107d;
	-- d109d
	sted109d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord109d,
			Enable=>Enabled109d,
			match=>matchd109d,
			run=>run);

	Enabled109d <= matchd109d OR matchd108d;
	-- d110d
	sted110d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord110d,
			Enable=>Enabled110d,
			match=>matchd110d,
			run=>run);

	reports(7) <= matchd110d;
	Enabled110d <= matchd109d;
	-- d111d
	sted111d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord111d,
			Enable=>Enabled111d,
			match=>matchd111d,
			run=>run);

	-- d112d
	sted112d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord112d,
			Enable=>Enabled112d,
			match=>matchd112d,
			run=>run);

	Enabled112d <= matchd112d OR matchd111d;
	-- d113d
	sted113d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord113d,
			Enable=>Enabled113d,
			match=>matchd113d,
			run=>run);

	Enabled113d <= matchd112d;
	-- d114d
	sted114d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord114d,
			Enable=>Enabled114d,
			match=>matchd114d,
			run=>run);

	Enabled114d <= matchd113d;
	-- d115d
	sted115d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord115d,
			Enable=>Enabled115d,
			match=>matchd115d,
			run=>run);

	Enabled115d <= matchd114d;
	-- d116d
	sted116d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord116d,
			Enable=>Enabled116d,
			match=>matchd116d,
			run=>run);

	Enabled116d <= matchd115d;
	-- d117d
	sted117d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord117d,
			Enable=>Enabled117d,
			match=>matchd117d,
			run=>run);

	Enabled117d <= matchd116d;
	-- d118d
	sted118d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord118d,
			Enable=>Enabled118d,
			match=>matchd118d,
			run=>run);

	Enabled118d <= matchd117d;
	-- d119d
	sted119d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord119d,
			Enable=>Enabled119d,
			match=>matchd119d,
			run=>run);

	Enabled119d <= matchd118d;
	-- d120d
	sted120d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord120d,
			Enable=>Enabled120d,
			match=>matchd120d,
			run=>run);

	Enabled120d <= matchd119d;
	-- d121d
	sted121d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord121d,
			Enable=>Enabled121d,
			match=>matchd121d,
			run=>run);

	Enabled121d <= matchd121d OR matchd120d;
	-- d122d
	sted122d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord122d,
			Enable=>Enabled122d,
			match=>matchd122d,
			run=>run);

	reports(8) <= matchd122d;
	Enabled122d <= matchd121d;
	-- d123d
	sted123d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord123d,
			Enable=>Enabled123d,
			match=>matchd123d,
			run=>run);

	-- d124d
	sted124d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord124d,
			Enable=>Enabled124d,
			match=>matchd124d,
			run=>run);

	Enabled124d <= matchd123d;
	-- d125d
	sted125d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord125d,
			Enable=>Enabled125d,
			match=>matchd125d,
			run=>run);

	Enabled125d <= matchd124d;
	-- d126d
	sted126d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord126d,
			Enable=>Enabled126d,
			match=>matchd126d,
			run=>run);

	Enabled126d <= matchd125d;
	-- d127d
	sted127d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord127d,
			Enable=>Enabled127d,
			match=>matchd127d,
			run=>run);

	Enabled127d <= matchd126d;
	-- d128d
	sted128d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord128d,
			Enable=>Enabled128d,
			match=>matchd128d,
			run=>run);

	Enabled128d <= matchd128d OR matchd127d;
	-- d129d
	sted129d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord129d,
			Enable=>Enabled129d,
			match=>matchd129d,
			run=>run);

	Enabled129d <= matchd128d;
	-- d130d
	sted130d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord130d,
			Enable=>Enabled130d,
			match=>matchd130d,
			run=>run);

	Enabled130d <= matchd129d;
	-- d131d
	sted131d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord131d,
			Enable=>Enabled131d,
			match=>matchd131d,
			run=>run);

	Enabled131d <= matchd130d;
	-- d132d
	sted132d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord132d,
			Enable=>Enabled132d,
			match=>matchd132d,
			run=>run);

	Enabled132d <= matchd131d;
	-- d133d
	sted133d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord133d,
			Enable=>Enabled133d,
			match=>matchd133d,
			run=>run);

	Enabled133d <= matchd132d;
	-- d134d
	sted134d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord134d,
			Enable=>Enabled134d,
			match=>matchd134d,
			run=>run);

	Enabled134d <= matchd133d;
	-- d135d
	sted135d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord135d,
			Enable=>Enabled135d,
			match=>matchd135d,
			run=>run);

	Enabled135d <= matchd134d;
	-- d136d
	sted136d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord136d,
			Enable=>Enabled136d,
			match=>matchd136d,
			run=>run);

	Enabled136d <= matchd135d;
	-- d137d
	sted137d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord137d,
			Enable=>Enabled137d,
			match=>matchd137d,
			run=>run);

	reports(9) <= matchd137d;
	Enabled137d <= matchd136d;
	-- d138d
	sted138d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord138d,
			Enable=>Enabled138d,
			match=>matchd138d,
			run=>run);

	-- d139d
	sted139d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord139d,
			Enable=>Enabled139d,
			match=>matchd139d,
			run=>run);

	Enabled139d <= matchd138d;
	-- d140d
	sted140d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord140d,
			Enable=>Enabled140d,
			match=>matchd140d,
			run=>run);

	Enabled140d <= matchd139d;
	-- d141d
	sted141d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord141d,
			Enable=>Enabled141d,
			match=>matchd141d,
			run=>run);

	Enabled141d <= matchd140d;
	-- d142d
	sted142d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord142d,
			Enable=>Enabled142d,
			match=>matchd142d,
			run=>run);

	Enabled142d <= matchd141d;
	-- d143d
	sted143d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord143d,
			Enable=>Enabled143d,
			match=>matchd143d,
			run=>run);

	Enabled143d <= matchd142d;
	-- d144d
	sted144d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord144d,
			Enable=>Enabled144d,
			match=>matchd144d,
			run=>run);

	Enabled144d <= matchd143d;
	-- d145d
	sted145d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord145d,
			Enable=>Enabled145d,
			match=>matchd145d,
			run=>run);

	Enabled145d <= matchd144d;
	-- d146d
	sted146d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord146d,
			Enable=>Enabled146d,
			match=>matchd146d,
			run=>run);

	Enabled146d <= matchd145d;
	-- d147d
	sted147d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord147d,
			Enable=>Enabled147d,
			match=>matchd147d,
			run=>run);

	Enabled147d <= matchd146d;
	-- d148d
	sted148d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord148d,
			Enable=>Enabled148d,
			match=>matchd148d,
			run=>run);

	Enabled148d <= matchd147d;
	-- d149d
	sted149d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord149d,
			Enable=>Enabled149d,
			match=>matchd149d,
			run=>run);

	Enabled149d <= matchd148d;
	-- d150d
	sted150d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord150d,
			Enable=>Enabled150d,
			match=>matchd150d,
			run=>run);

	Enabled150d <= matchd150d OR matchd149d;
	-- d151d
	sted151d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord151d,
			Enable=>Enabled151d,
			match=>matchd151d,
			run=>run);

	reports(10) <= matchd151d;
	Enabled151d <= matchd150d;
	-- d152d
	sted152d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord152d,
			Enable=>Enabled152d,
			match=>matchd152d,
			run=>run);

	-- d153d
	sted153d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord153d,
			Enable=>Enabled153d,
			match=>matchd153d,
			run=>run);

	Enabled153d <= matchd152d OR matchd153d;
	-- d154d
	sted154d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord154d,
			Enable=>Enabled154d,
			match=>matchd154d,
			run=>run);

	Enabled154d <= matchd153d;
	-- d155d
	sted155d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord155d,
			Enable=>Enabled155d,
			match=>matchd155d,
			run=>run);

	Enabled155d <= matchd154d;
	-- d156d
	sted156d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord156d,
			Enable=>Enabled156d,
			match=>matchd156d,
			run=>run);

	Enabled156d <= matchd155d;
	-- d157d
	sted157d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord157d,
			Enable=>Enabled157d,
			match=>matchd157d,
			run=>run);

	Enabled157d <= matchd156d;
	-- d158d
	sted158d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord158d,
			Enable=>Enabled158d,
			match=>matchd158d,
			run=>run);

	Enabled158d <= matchd157d;
	-- d159d
	sted159d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord159d,
			Enable=>Enabled159d,
			match=>matchd159d,
			run=>run);

	Enabled159d <= matchd158d;
	-- d160d
	sted160d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord160d,
			Enable=>Enabled160d,
			match=>matchd160d,
			run=>run);

	Enabled160d <= matchd159d;
	-- d161d
	sted161d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord161d,
			Enable=>Enabled161d,
			match=>matchd161d,
			run=>run);

	Enabled161d <= matchd160d;
	-- d162d
	sted162d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord162d,
			Enable=>Enabled162d,
			match=>matchd162d,
			run=>run);

	Enabled162d <= matchd161d;
	-- d163d
	sted163d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord163d,
			Enable=>Enabled163d,
			match=>matchd163d,
			run=>run);

	Enabled163d <= matchd162d;
	-- d164d
	sted164d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord164d,
			Enable=>Enabled164d,
			match=>matchd164d,
			run=>run);

	Enabled164d <= matchd164d OR matchd163d;
	-- d165d
	sted165d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord165d,
			Enable=>Enabled165d,
			match=>matchd165d,
			run=>run);

	reports(11) <= matchd165d;
	Enabled165d <= matchd164d;
	-- d166d
	sted166d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord166d,
			Enable=>Enabled166d,
			match=>matchd166d,
			run=>run);

	-- d167d
	sted167d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord167d,
			Enable=>Enabled167d,
			match=>matchd167d,
			run=>run);

	Enabled167d <= matchd167d OR matchd166d;
	-- d168d
	sted168d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord168d,
			Enable=>Enabled168d,
			match=>matchd168d,
			run=>run);

	Enabled168d <= matchd167d;
	-- d169d
	sted169d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord169d,
			Enable=>Enabled169d,
			match=>matchd169d,
			run=>run);

	Enabled169d <= matchd168d;
	-- d170d
	sted170d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord170d,
			Enable=>Enabled170d,
			match=>matchd170d,
			run=>run);

	Enabled170d <= matchd169d;
	-- d171d
	sted171d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord171d,
			Enable=>Enabled171d,
			match=>matchd171d,
			run=>run);

	Enabled171d <= matchd170d;
	-- d172d
	sted172d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord172d,
			Enable=>Enabled172d,
			match=>matchd172d,
			run=>run);

	Enabled172d <= matchd171d;
	-- d173d
	sted173d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord173d,
			Enable=>Enabled173d,
			match=>matchd173d,
			run=>run);

	Enabled173d <= matchd172d;
	-- d174d
	sted174d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord174d,
			Enable=>Enabled174d,
			match=>matchd174d,
			run=>run);

	Enabled174d <= matchd173d;
	-- d175d
	sted175d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord175d,
			Enable=>Enabled175d,
			match=>matchd175d,
			run=>run);

	Enabled175d <= matchd174d OR matchd175d;
	-- d176d
	sted176d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord176d,
			Enable=>Enabled176d,
			match=>matchd176d,
			run=>run);

	reports(12) <= matchd176d;
	Enabled176d <= matchd175d;
	-- d177d
	sted177d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord177d,
			Enable=>Enabled177d,
			match=>matchd177d,
			run=>run);

	-- d178d
	sted178d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord178d,
			Enable=>Enabled178d,
			match=>matchd178d,
			run=>run);

	Enabled178d <= matchd177d OR matchd178d;
	-- d179d
	sted179d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord179d,
			Enable=>Enabled179d,
			match=>matchd179d,
			run=>run);

	Enabled179d <= matchd178d;
	-- d180d
	sted180d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord180d,
			Enable=>Enabled180d,
			match=>matchd180d,
			run=>run);

	Enabled180d <= matchd179d;
	-- d181d
	sted181d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord181d,
			Enable=>Enabled181d,
			match=>matchd181d,
			run=>run);

	Enabled181d <= matchd180d;
	-- d182d
	sted182d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord182d,
			Enable=>Enabled182d,
			match=>matchd182d,
			run=>run);

	Enabled182d <= matchd181d;
	-- d183d
	sted183d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord183d,
			Enable=>Enabled183d,
			match=>matchd183d,
			run=>run);

	Enabled183d <= matchd182d;
	-- d184d
	sted184d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord184d,
			Enable=>Enabled184d,
			match=>matchd184d,
			run=>run);

	Enabled184d <= matchd183d;
	-- d185d
	sted185d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord185d,
			Enable=>Enabled185d,
			match=>matchd185d,
			run=>run);

	Enabled185d <= matchd184d;
	-- d186d
	sted186d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord186d,
			Enable=>Enabled186d,
			match=>matchd186d,
			run=>run);

	Enabled186d <= matchd185d OR matchd186d;
	-- d187d
	sted187d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord187d,
			Enable=>Enabled187d,
			match=>matchd187d,
			run=>run);

	reports(13) <= matchd187d;
	Enabled187d <= matchd186d;
	-- d188d
	sted188d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord188d,
			Enable=>Enabled188d,
			match=>matchd188d,
			run=>run);

	-- d189d
	sted189d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord189d,
			Enable=>Enabled189d,
			match=>matchd189d,
			run=>run);

	Enabled189d <= matchd188d;
	-- d190d
	sted190d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord190d,
			Enable=>Enabled190d,
			match=>matchd190d,
			run=>run);

	Enabled190d <= matchd189d;
	-- d191d
	sted191d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord191d,
			Enable=>Enabled191d,
			match=>matchd191d,
			run=>run);

	Enabled191d <= matchd190d;
	-- d192d
	sted192d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord192d,
			Enable=>Enabled192d,
			match=>matchd192d,
			run=>run);

	Enabled192d <= matchd191d;
	-- d193d
	sted193d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord193d,
			Enable=>Enabled193d,
			match=>matchd193d,
			run=>run);

	Enabled193d <= matchd192d;
	-- d194d
	sted194d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord194d,
			Enable=>Enabled194d,
			match=>matchd194d,
			run=>run);

	Enabled194d <= matchd193d;
	-- d195d
	sted195d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord195d,
			Enable=>Enabled195d,
			match=>matchd195d,
			run=>run);

	Enabled195d <= matchd194d;
	-- d196d
	sted196d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord196d,
			Enable=>Enabled196d,
			match=>matchd196d,
			run=>run);

	Enabled196d <= matchd195d;
	-- d197d
	sted197d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord197d,
			Enable=>Enabled197d,
			match=>matchd197d,
			run=>run);

	Enabled197d <= matchd196d;
	-- d198d
	sted198d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord198d,
			Enable=>Enabled198d,
			match=>matchd198d,
			run=>run);

	Enabled198d <= matchd197d;
	-- d199d
	sted199d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord199d,
			Enable=>Enabled199d,
			match=>matchd199d,
			run=>run);

	Enabled199d <= matchd198d OR matchd199d;
	-- d200d
	sted200d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord200d,
			Enable=>Enabled200d,
			match=>matchd200d,
			run=>run);

	reports(14) <= matchd200d;
	Enabled200d <= matchd199d;
	-- d201d
	sted201d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord201d,
			Enable=>Enabled201d,
			match=>matchd201d,
			run=>run);

	-- d202d
	sted202d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord202d,
			Enable=>Enabled202d,
			match=>matchd202d,
			run=>run);

	Enabled202d <= matchd201d;
	-- d203d
	sted203d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord203d,
			Enable=>Enabled203d,
			match=>matchd203d,
			run=>run);

	Enabled203d <= matchd202d;
	-- d204d
	sted204d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord204d,
			Enable=>Enabled204d,
			match=>matchd204d,
			run=>run);

	Enabled204d <= matchd203d;
	-- d205d
	sted205d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord205d,
			Enable=>Enabled205d,
			match=>matchd205d,
			run=>run);

	Enabled205d <= matchd204d;
	-- d206d
	sted206d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord206d,
			Enable=>Enabled206d,
			match=>matchd206d,
			run=>run);

	Enabled206d <= matchd205d;
	-- d207d
	sted207d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord207d,
			Enable=>Enabled207d,
			match=>matchd207d,
			run=>run);

	Enabled207d <= matchd206d;
	-- d208d
	sted208d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord208d,
			Enable=>Enabled208d,
			match=>matchd208d,
			run=>run);

	Enabled208d <= matchd207d;
	-- d209d
	sted209d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord209d,
			Enable=>Enabled209d,
			match=>matchd209d,
			run=>run);

	Enabled209d <= matchd208d;
	-- d210d
	sted210d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord210d,
			Enable=>Enabled210d,
			match=>matchd210d,
			run=>run);

	Enabled210d <= matchd209d OR matchd210d;
	-- d211d
	sted211d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord211d,
			Enable=>Enabled211d,
			match=>matchd211d,
			run=>run);

	reports(15) <= matchd211d;
	Enabled211d <= matchd210d;
	-- d212d
	sted212d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord212d,
			Enable=>Enabled212d,
			match=>matchd212d,
			run=>run);

	-- d213d
	sted213d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord213d,
			Enable=>Enabled213d,
			match=>matchd213d,
			run=>run);

	Enabled213d <= matchd213d OR matchd212d;
	-- d214d
	sted214d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord214d,
			Enable=>Enabled214d,
			match=>matchd214d,
			run=>run);

	Enabled214d <= matchd213d;
	-- d215d
	sted215d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord215d,
			Enable=>Enabled215d,
			match=>matchd215d,
			run=>run);

	Enabled215d <= matchd214d;
	-- d216d
	sted216d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord216d,
			Enable=>Enabled216d,
			match=>matchd216d,
			run=>run);

	Enabled216d <= matchd215d;
	-- d217d
	sted217d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord217d,
			Enable=>Enabled217d,
			match=>matchd217d,
			run=>run);

	Enabled217d <= matchd216d;
	-- d218d
	sted218d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord218d,
			Enable=>Enabled218d,
			match=>matchd218d,
			run=>run);

	Enabled218d <= matchd218d OR matchd217d;
	-- d219d
	sted219d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord219d,
			Enable=>Enabled219d,
			match=>matchd219d,
			run=>run);

	Enabled219d <= matchd218d;
	-- d220d
	sted220d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord220d,
			Enable=>Enabled220d,
			match=>matchd220d,
			run=>run);

	Enabled220d <= matchd219d;
	-- d221d
	sted221d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord221d,
			Enable=>Enabled221d,
			match=>matchd221d,
			run=>run);

	Enabled221d <= matchd220d;
	-- d222d
	sted222d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord222d,
			Enable=>Enabled222d,
			match=>matchd222d,
			run=>run);

	reports(16) <= matchd222d;
	Enabled222d <= matchd221d;
	-- d223d
	sted223d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord223d,
			Enable=>Enabled223d,
			match=>matchd223d,
			run=>run);

	-- d224d
	sted224d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord224d,
			Enable=>Enabled224d,
			match=>matchd224d,
			run=>run);

	Enabled224d <= matchd223d OR matchd224d;
	-- d225d
	sted225d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord225d,
			Enable=>Enabled225d,
			match=>matchd225d,
			run=>run);

	Enabled225d <= matchd224d;
	-- d226d
	sted226d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord226d,
			Enable=>Enabled226d,
			match=>matchd226d,
			run=>run);

	Enabled226d <= matchd225d;
	-- d227d
	sted227d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord227d,
			Enable=>Enabled227d,
			match=>matchd227d,
			run=>run);

	Enabled227d <= matchd226d;
	-- d228d
	sted228d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord228d,
			Enable=>Enabled228d,
			match=>matchd228d,
			run=>run);

	Enabled228d <= matchd227d;
	-- d229d
	sted229d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord229d,
			Enable=>Enabled229d,
			match=>matchd229d,
			run=>run);

	Enabled229d <= matchd228d;
	-- d230d
	sted230d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord230d,
			Enable=>Enabled230d,
			match=>matchd230d,
			run=>run);

	Enabled230d <= matchd229d OR matchd230d;
	-- d231d
	sted231d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord231d,
			Enable=>Enabled231d,
			match=>matchd231d,
			run=>run);

	Enabled231d <= matchd230d;
	-- d232d
	sted232d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord232d,
			Enable=>Enabled232d,
			match=>matchd232d,
			run=>run);

	Enabled232d <= matchd231d;
	-- d233d
	sted233d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord233d,
			Enable=>Enabled233d,
			match=>matchd233d,
			run=>run);

	Enabled233d <= matchd232d;
	-- d234d
	sted234d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord234d,
			Enable=>Enabled234d,
			match=>matchd234d,
			run=>run);

	reports(17) <= matchd234d;
	Enabled234d <= matchd233d;
	-- d235d
	sted235d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord235d,
			Enable=>Enabled235d,
			match=>matchd235d,
			run=>run);

	-- d236d
	sted236d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord236d,
			Enable=>Enabled236d,
			match=>matchd236d,
			run=>run);

	Enabled236d <= matchd236d OR matchd235d;
	-- d237d
	sted237d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord237d,
			Enable=>Enabled237d,
			match=>matchd237d,
			run=>run);

	Enabled237d <= matchd236d;
	-- d238d
	sted238d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord238d,
			Enable=>Enabled238d,
			match=>matchd238d,
			run=>run);

	Enabled238d <= matchd238d OR matchd237d;
	-- d239d
	sted239d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord239d,
			Enable=>Enabled239d,
			match=>matchd239d,
			run=>run);

	Enabled239d <= matchd238d;
	-- d240d
	sted240d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord240d,
			Enable=>Enabled240d,
			match=>matchd240d,
			run=>run);

	Enabled240d <= matchd239d OR matchd240d;
	-- d241d
	sted241d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord241d,
			Enable=>Enabled241d,
			match=>matchd241d,
			run=>run);

	Enabled241d <= matchd240d;
	-- d242d
	sted242d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord242d,
			Enable=>Enabled242d,
			match=>matchd242d,
			run=>run);

	Enabled242d <= matchd241d;
	-- d243d
	sted243d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord243d,
			Enable=>Enabled243d,
			match=>matchd243d,
			run=>run);

	Enabled243d <= matchd242d;
	-- d244d
	sted244d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord244d,
			Enable=>Enabled244d,
			match=>matchd244d,
			run=>run);

	Enabled244d <= matchd243d;
	-- d245d
	sted245d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord245d,
			Enable=>Enabled245d,
			match=>matchd245d,
			run=>run);

	Enabled245d <= matchd244d;
	-- d246d
	sted246d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord246d,
			Enable=>Enabled246d,
			match=>matchd246d,
			run=>run);

	Enabled246d <= matchd246d OR matchd245d;
	-- d247d
	sted247d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord247d,
			Enable=>Enabled247d,
			match=>matchd247d,
			run=>run);

	Enabled247d <= matchd246d;
	-- d248d
	sted248d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord248d,
			Enable=>Enabled248d,
			match=>matchd248d,
			run=>run);

	Enabled248d <= matchd247d;
	-- d249d
	sted249d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord249d,
			Enable=>Enabled249d,
			match=>matchd249d,
			run=>run);

	Enabled249d <= matchd248d;
	-- d250d
	sted250d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord250d,
			Enable=>Enabled250d,
			match=>matchd250d,
			run=>run);

	Enabled250d <= matchd249d;
	-- d251d
	sted251d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord251d,
			Enable=>Enabled251d,
			match=>matchd251d,
			run=>run);

	Enabled251d <= matchd250d;
	-- d252d
	sted252d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord252d,
			Enable=>Enabled252d,
			match=>matchd252d,
			run=>run);

	-- d253d
	sted253d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord253d,
			Enable=>Enabled253d,
			match=>matchd253d,
			run=>run);

	Enabled253d <= matchd253d OR matchd252d;
	-- d254d
	sted254d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord254d,
			Enable=>Enabled254d,
			match=>matchd254d,
			run=>run);

	Enabled254d <= matchd253d;
	-- d255d
	sted255d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord255d,
			Enable=>Enabled255d,
			match=>matchd255d,
			run=>run);

	Enabled255d <= matchd254d;
	-- d256d
	sted256d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord256d,
			Enable=>Enabled256d,
			match=>matchd256d,
			run=>run);

	Enabled256d <= matchd255d;
	-- d257d
	sted257d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord257d,
			Enable=>Enabled257d,
			match=>matchd257d,
			run=>run);

	Enabled257d <= matchd256d;
	-- d258d
	sted258d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord258d,
			Enable=>Enabled258d,
			match=>matchd258d,
			run=>run);

	Enabled258d <= matchd257d;
	-- d259d
	sted259d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord259d,
			Enable=>Enabled259d,
			match=>matchd259d,
			run=>run);

	Enabled259d <= matchd259d OR matchd258d;
	-- d260d
	sted260d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord260d,
			Enable=>Enabled260d,
			match=>matchd260d,
			run=>run);

	Enabled260d <= matchd259d;
	-- d261d
	sted261d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord261d,
			Enable=>Enabled261d,
			match=>matchd261d,
			run=>run);

	Enabled261d <= matchd260d OR matchd261d;
	-- d262d
	sted262d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord262d,
			Enable=>Enabled262d,
			match=>matchd262d,
			run=>run);

	Enabled262d <= matchd261d;
	-- d263d
	sted263d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord263d,
			Enable=>Enabled263d,
			match=>matchd263d,
			run=>run);

	Enabled263d <= matchd262d OR matchd263d;
	-- d264d
	sted264d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord264d,
			Enable=>Enabled264d,
			match=>matchd264d,
			run=>run);

	Enabled264d <= matchd263d;
	-- d265d
	sted265d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord265d,
			Enable=>Enabled265d,
			match=>matchd265d,
			run=>run);

	Enabled265d <= matchd264d;
	-- d266d
	sted266d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord266d,
			Enable=>Enabled266d,
			match=>matchd266d,
			run=>run);

	Enabled266d <= matchd265d;
	-- d267d
	sted267d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord267d,
			Enable=>Enabled267d,
			match=>matchd267d,
			run=>run);

	Enabled267d <= matchd266d;
	-- d268d
	sted268d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord268d,
			Enable=>Enabled268d,
			match=>matchd268d,
			run=>run);

	Enabled268d <= matchd267d;
	-- d270d
	sted270d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord270d,
			Enable=>Enabled270d,
			match=>matchd270d,
			run=>run);

	-- d271d
	sted271d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord271d,
			Enable=>Enabled271d,
			match=>matchd271d,
			run=>run);

	Enabled271d <= matchd271d OR matchd270d;
	-- d272d
	sted272d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord272d,
			Enable=>Enabled272d,
			match=>matchd272d,
			run=>run);

	Enabled272d <= matchd271d;
	-- d273d
	sted273d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord273d,
			Enable=>Enabled273d,
			match=>matchd273d,
			run=>run);

	Enabled273d <= matchd272d;
	-- d274d
	sted274d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord274d,
			Enable=>Enabled274d,
			match=>matchd274d,
			run=>run);

	Enabled274d <= matchd273d;
	-- d275d
	sted275d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord275d,
			Enable=>Enabled275d,
			match=>matchd275d,
			run=>run);

	Enabled275d <= matchd274d;
	-- d276d
	sted276d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord276d,
			Enable=>Enabled276d,
			match=>matchd276d,
			run=>run);

	Enabled276d <= matchd275d;
	-- d277d
	sted277d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord277d,
			Enable=>Enabled277d,
			match=>matchd277d,
			run=>run);

	Enabled277d <= matchd277d OR matchd276d;
	-- d278d
	sted278d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord278d,
			Enable=>Enabled278d,
			match=>matchd278d,
			run=>run);

	Enabled278d <= matchd277d;
	-- d279d
	sted279d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord279d,
			Enable=>Enabled279d,
			match=>matchd279d,
			run=>run);

	Enabled279d <= matchd278d;
	-- d280d
	sted280d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord280d,
			Enable=>Enabled280d,
			match=>matchd280d,
			run=>run);

	Enabled280d <= matchd279d;
	-- d281d
	sted281d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord281d,
			Enable=>Enabled281d,
			match=>matchd281d,
			run=>run);

	Enabled281d <= matchd280d;
	-- d282d
	sted282d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord282d,
			Enable=>Enabled282d,
			match=>matchd282d,
			run=>run);

	reports(18) <= matchd282d;
	Enabled282d <= matchd281d;
	-- d283d
	sted283d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord283d,
			Enable=>Enabled283d,
			match=>matchd283d,
			run=>run);

	-- d284d
	sted284d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord284d,
			Enable=>Enabled284d,
			match=>matchd284d,
			run=>run);

	Enabled284d <= matchd284d OR matchd283d;
	-- d285d
	sted285d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord285d,
			Enable=>Enabled285d,
			match=>matchd285d,
			run=>run);

	Enabled285d <= matchd284d;
	-- d286d
	sted286d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord286d,
			Enable=>Enabled286d,
			match=>matchd286d,
			run=>run);

	Enabled286d <= matchd286d OR matchd285d;
	-- d287d
	sted287d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord287d,
			Enable=>Enabled287d,
			match=>matchd287d,
			run=>run);

	Enabled287d <= matchd286d;
	-- d288d
	sted288d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord288d,
			Enable=>Enabled288d,
			match=>matchd288d,
			run=>run);

	Enabled288d <= matchd288d OR matchd287d;
	-- d289d
	sted289d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord289d,
			Enable=>Enabled289d,
			match=>matchd289d,
			run=>run);

	Enabled289d <= matchd288d;
	-- d290d
	sted290d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord290d,
			Enable=>Enabled290d,
			match=>matchd290d,
			run=>run);

	Enabled290d <= matchd289d;
	-- d291d
	sted291d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord291d,
			Enable=>Enabled291d,
			match=>matchd291d,
			run=>run);

	Enabled291d <= matchd290d;
	-- d292d
	sted292d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord292d,
			Enable=>Enabled292d,
			match=>matchd292d,
			run=>run);

	Enabled292d <= matchd291d;
	-- d293d
	sted293d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord293d,
			Enable=>Enabled293d,
			match=>matchd293d,
			run=>run);

	Enabled293d <= matchd293d OR matchd292d;
	-- d294d
	sted294d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord294d,
			Enable=>Enabled294d,
			match=>matchd294d,
			run=>run);

	Enabled294d <= matchd293d;
	-- d295d
	sted295d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord295d,
			Enable=>Enabled295d,
			match=>matchd295d,
			run=>run);

	Enabled295d <= matchd294d;
	-- d296d
	sted296d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord296d,
			Enable=>Enabled296d,
			match=>matchd296d,
			run=>run);

	Enabled296d <= matchd295d;
	-- d297d
	sted297d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord297d,
			Enable=>Enabled297d,
			match=>matchd297d,
			run=>run);

	Enabled297d <= matchd296d;
	-- d298d
	sted298d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord298d,
			Enable=>Enabled298d,
			match=>matchd298d,
			run=>run);

	-- d299d
	sted299d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord299d,
			Enable=>Enabled299d,
			match=>matchd299d,
			run=>run);

	Enabled299d <= matchd298d OR matchd299d;
	-- d300d
	sted300d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord300d,
			Enable=>Enabled300d,
			match=>matchd300d,
			run=>run);

	Enabled300d <= matchd299d;
	-- d301d
	sted301d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord301d,
			Enable=>Enabled301d,
			match=>matchd301d,
			run=>run);

	Enabled301d <= matchd300d;
	-- d302d
	sted302d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord302d,
			Enable=>Enabled302d,
			match=>matchd302d,
			run=>run);

	Enabled302d <= matchd301d;
	-- d303d
	sted303d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord303d,
			Enable=>Enabled303d,
			match=>matchd303d,
			run=>run);

	Enabled303d <= matchd302d;
	-- d304d
	sted304d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord304d,
			Enable=>Enabled304d,
			match=>matchd304d,
			run=>run);

	Enabled304d <= matchd304d OR matchd303d;
	-- d305d
	sted305d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord305d,
			Enable=>Enabled305d,
			match=>matchd305d,
			run=>run);

	Enabled305d <= matchd304d;
	-- d306d
	sted306d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord306d,
			Enable=>Enabled306d,
			match=>matchd306d,
			run=>run);

	Enabled306d <= matchd306d OR matchd305d;
	-- d307d
	sted307d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord307d,
			Enable=>Enabled307d,
			match=>matchd307d,
			run=>run);

	Enabled307d <= matchd306d;
	-- d308d
	sted308d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord308d,
			Enable=>Enabled308d,
			match=>matchd308d,
			run=>run);

	Enabled308d <= matchd307d OR matchd308d;
	-- d309d
	sted309d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord309d,
			Enable=>Enabled309d,
			match=>matchd309d,
			run=>run);

	Enabled309d <= matchd308d;
	-- d310d
	sted310d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord310d,
			Enable=>Enabled310d,
			match=>matchd310d,
			run=>run);

	Enabled310d <= matchd309d;
	-- d311d
	sted311d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord311d,
			Enable=>Enabled311d,
			match=>matchd311d,
			run=>run);

	Enabled311d <= matchd310d;
	-- d312d
	sted312d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord312d,
			Enable=>Enabled312d,
			match=>matchd312d,
			run=>run);

	Enabled312d <= matchd311d;
	-- d314d
	sted314d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord314d,
			Enable=>Enabled314d,
			match=>matchd314d,
			run=>run);

	-- d315d
	sted315d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord315d,
			Enable=>Enabled315d,
			match=>matchd315d,
			run=>run);

	Enabled315d <= matchd315d OR matchd314d;
	-- d316d
	sted316d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord316d,
			Enable=>Enabled316d,
			match=>matchd316d,
			run=>run);

	Enabled316d <= matchd315d;
	-- d317d
	sted317d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord317d,
			Enable=>Enabled317d,
			match=>matchd317d,
			run=>run);

	Enabled317d <= matchd316d;
	-- d318d
	sted318d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord318d,
			Enable=>Enabled318d,
			match=>matchd318d,
			run=>run);

	Enabled318d <= matchd317d;
	-- d319d
	sted319d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord319d,
			Enable=>Enabled319d,
			match=>matchd319d,
			run=>run);

	Enabled319d <= matchd318d;
	-- d320d
	sted320d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord320d,
			Enable=>Enabled320d,
			match=>matchd320d,
			run=>run);

	Enabled320d <= matchd319d;
	-- d321d
	sted321d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord321d,
			Enable=>Enabled321d,
			match=>matchd321d,
			run=>run);

	Enabled321d <= matchd321d OR matchd320d;
	-- d322d
	sted322d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord322d,
			Enable=>Enabled322d,
			match=>matchd322d,
			run=>run);

	Enabled322d <= matchd321d;
	-- d323d
	sted323d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord323d,
			Enable=>Enabled323d,
			match=>matchd323d,
			run=>run);

	Enabled323d <= matchd322d;
	-- d324d
	sted324d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord324d,
			Enable=>Enabled324d,
			match=>matchd324d,
			run=>run);

	Enabled324d <= matchd323d;
	-- d325d
	sted325d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord325d,
			Enable=>Enabled325d,
			match=>matchd325d,
			run=>run);

	reports(19) <= matchd325d;
	Enabled325d <= matchd324d;
	-- d326d
	sted326d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord326d,
			Enable=>Enabled326d,
			match=>matchd326d,
			run=>run);

	-- d327d
	sted327d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord327d,
			Enable=>Enabled327d,
			match=>matchd327d,
			run=>run);

	Enabled327d <= matchd327d OR matchd326d;
	-- d328d
	sted328d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord328d,
			Enable=>Enabled328d,
			match=>matchd328d,
			run=>run);

	Enabled328d <= matchd327d;
	-- d329d
	sted329d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord329d,
			Enable=>Enabled329d,
			match=>matchd329d,
			run=>run);

	Enabled329d <= matchd329d OR matchd328d;
	-- d330d
	sted330d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord330d,
			Enable=>Enabled330d,
			match=>matchd330d,
			run=>run);

	Enabled330d <= matchd329d;
	-- d331d
	sted331d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord331d,
			Enable=>Enabled331d,
			match=>matchd331d,
			run=>run);

	Enabled331d <= matchd330d OR matchd331d;
	-- d332d
	sted332d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord332d,
			Enable=>Enabled332d,
			match=>matchd332d,
			run=>run);

	Enabled332d <= matchd331d;
	-- d333d
	sted333d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord333d,
			Enable=>Enabled333d,
			match=>matchd333d,
			run=>run);

	Enabled333d <= matchd332d;
	-- d334d
	sted334d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord334d,
			Enable=>Enabled334d,
			match=>matchd334d,
			run=>run);

	Enabled334d <= matchd333d;
	-- d335d
	sted335d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord335d,
			Enable=>Enabled335d,
			match=>matchd335d,
			run=>run);

	Enabled335d <= matchd334d;
	-- d336d
	sted336d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord336d,
			Enable=>Enabled336d,
			match=>matchd336d,
			run=>run);

	Enabled336d <= matchd336d OR matchd335d;
	-- d337d
	sted337d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord337d,
			Enable=>Enabled337d,
			match=>matchd337d,
			run=>run);

	Enabled337d <= matchd336d;
	-- d338d
	sted338d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord338d,
			Enable=>Enabled338d,
			match=>matchd338d,
			run=>run);

	Enabled338d <= matchd337d;
	-- d339d
	sted339d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord339d,
			Enable=>Enabled339d,
			match=>matchd339d,
			run=>run);

	Enabled339d <= matchd338d;
	-- d340d
	sted340d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord340d,
			Enable=>Enabled340d,
			match=>matchd340d,
			run=>run);

	Enabled340d <= matchd339d;
	-- d341d
	sted341d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord341d,
			Enable=>Enabled341d,
			match=>matchd341d,
			run=>run);

	-- d342d
	sted342d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord342d,
			Enable=>Enabled342d,
			match=>matchd342d,
			run=>run);

	Enabled342d <= matchd342d OR matchd341d;
	-- d343d
	sted343d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord343d,
			Enable=>Enabled343d,
			match=>matchd343d,
			run=>run);

	Enabled343d <= matchd342d;
	-- d344d
	sted344d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord344d,
			Enable=>Enabled344d,
			match=>matchd344d,
			run=>run);

	Enabled344d <= matchd343d;
	-- d345d
	sted345d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord345d,
			Enable=>Enabled345d,
			match=>matchd345d,
			run=>run);

	Enabled345d <= matchd344d;
	-- d346d
	sted346d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord346d,
			Enable=>Enabled346d,
			match=>matchd346d,
			run=>run);

	Enabled346d <= matchd345d;
	-- d347d
	sted347d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord347d,
			Enable=>Enabled347d,
			match=>matchd347d,
			run=>run);

	Enabled347d <= matchd347d OR matchd346d;
	-- d348d
	sted348d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord348d,
			Enable=>Enabled348d,
			match=>matchd348d,
			run=>run);

	Enabled348d <= matchd347d;
	-- d349d
	sted349d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord349d,
			Enable=>Enabled349d,
			match=>matchd349d,
			run=>run);

	Enabled349d <= matchd349d OR matchd348d;
	-- d350d
	sted350d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord350d,
			Enable=>Enabled350d,
			match=>matchd350d,
			run=>run);

	Enabled350d <= matchd349d;
	-- d351d
	sted351d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord351d,
			Enable=>Enabled351d,
			match=>matchd351d,
			run=>run);

	Enabled351d <= matchd351d OR matchd350d;
	-- d352d
	sted352d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord352d,
			Enable=>Enabled352d,
			match=>matchd352d,
			run=>run);

	Enabled352d <= matchd351d;
	-- d353d
	sted353d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord353d,
			Enable=>Enabled353d,
			match=>matchd353d,
			run=>run);

	Enabled353d <= matchd352d;
	-- d354d
	sted354d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord354d,
			Enable=>Enabled354d,
			match=>matchd354d,
			run=>run);

	Enabled354d <= matchd353d;
	-- d355d
	sted355d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord355d,
			Enable=>Enabled355d,
			match=>matchd355d,
			run=>run);

	Enabled355d <= matchd354d;
	-- d357d
	sted357d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord357d,
			Enable=>Enabled357d,
			match=>matchd357d,
			run=>run);

	-- d358d
	sted358d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord358d,
			Enable=>Enabled358d,
			match=>matchd358d,
			run=>run);

	Enabled358d <= matchd358d OR matchd357d;
	-- d359d
	sted359d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord359d,
			Enable=>Enabled359d,
			match=>matchd359d,
			run=>run);

	Enabled359d <= matchd358d;
	-- d360d
	sted360d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord360d,
			Enable=>Enabled360d,
			match=>matchd360d,
			run=>run);

	Enabled360d <= matchd359d;
	-- d361d
	sted361d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord361d,
			Enable=>Enabled361d,
			match=>matchd361d,
			run=>run);

	Enabled361d <= matchd360d;
	-- d362d
	sted362d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord362d,
			Enable=>Enabled362d,
			match=>matchd362d,
			run=>run);

	Enabled362d <= matchd361d;
	-- d363d
	sted363d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord363d,
			Enable=>Enabled363d,
			match=>matchd363d,
			run=>run);

	Enabled363d <= matchd362d;
	-- d364d
	sted364d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord364d,
			Enable=>Enabled364d,
			match=>matchd364d,
			run=>run);

	Enabled364d <= matchd363d OR matchd364d;
	-- d365d
	sted365d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord365d,
			Enable=>Enabled365d,
			match=>matchd365d,
			run=>run);

	Enabled365d <= matchd364d;
	-- d366d
	sted366d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord366d,
			Enable=>Enabled366d,
			match=>matchd366d,
			run=>run);

	Enabled366d <= matchd365d;
	-- d367d
	sted367d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord367d,
			Enable=>Enabled367d,
			match=>matchd367d,
			run=>run);

	Enabled367d <= matchd366d;
	-- d368d
	sted368d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord368d,
			Enable=>Enabled368d,
			match=>matchd368d,
			run=>run);

	Enabled368d <= matchd367d;
	-- d369d
	sted369d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord369d,
			Enable=>Enabled369d,
			match=>matchd369d,
			run=>run);

	reports(20) <= matchd369d;
	Enabled369d <= matchd368d;
	-- d370d
	sted370d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord370d,
			Enable=>Enabled370d,
			match=>matchd370d,
			run=>run);

	-- d371d
	sted371d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord371d,
			Enable=>Enabled371d,
			match=>matchd371d,
			run=>run);

	Enabled371d <= matchd371d OR matchd370d;
	-- d372d
	sted372d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord372d,
			Enable=>Enabled372d,
			match=>matchd372d,
			run=>run);

	Enabled372d <= matchd371d;
	-- d373d
	sted373d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord373d,
			Enable=>Enabled373d,
			match=>matchd373d,
			run=>run);

	Enabled373d <= matchd372d;
	-- d374d
	sted374d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord374d,
			Enable=>Enabled374d,
			match=>matchd374d,
			run=>run);

	Enabled374d <= matchd373d;
	-- d375d
	sted375d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord375d,
			Enable=>Enabled375d,
			match=>matchd375d,
			run=>run);

	Enabled375d <= matchd374d;
	-- d376d
	sted376d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord376d,
			Enable=>Enabled376d,
			match=>matchd376d,
			run=>run);

	Enabled376d <= matchd375d;
	-- d377d
	sted377d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord377d,
			Enable=>Enabled377d,
			match=>matchd377d,
			run=>run);

	Enabled377d <= matchd376d OR matchd377d;
	-- d378d
	sted378d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord378d,
			Enable=>Enabled378d,
			match=>matchd378d,
			run=>run);

	Enabled378d <= matchd377d;
	-- d379d
	sted379d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord379d,
			Enable=>Enabled379d,
			match=>matchd379d,
			run=>run);

	Enabled379d <= matchd378d OR matchd379d;
	-- d380d
	sted380d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord380d,
			Enable=>Enabled380d,
			match=>matchd380d,
			run=>run);

	Enabled380d <= matchd379d;
	-- d381d
	sted381d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord381d,
			Enable=>Enabled381d,
			match=>matchd381d,
			run=>run);

	Enabled381d <= matchd381d OR matchd380d;
	-- d382d
	sted382d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord382d,
			Enable=>Enabled382d,
			match=>matchd382d,
			run=>run);

	Enabled382d <= matchd381d;
	-- d383d
	sted383d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord383d,
			Enable=>Enabled383d,
			match=>matchd383d,
			run=>run);

	Enabled383d <= matchd383d OR matchd382d;
	-- d384d
	sted384d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord384d,
			Enable=>Enabled384d,
			match=>matchd384d,
			run=>run);

	Enabled384d <= matchd383d;
	-- d385d
	sted385d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord385d,
			Enable=>Enabled385d,
			match=>matchd385d,
			run=>run);

	Enabled385d <= matchd385d OR matchd384d;
	-- d386d
	sted386d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord386d,
			Enable=>Enabled386d,
			match=>matchd386d,
			run=>run);

	Enabled386d <= matchd385d;
	-- d387d
	sted387d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord387d,
			Enable=>Enabled387d,
			match=>matchd387d,
			run=>run);

	Enabled387d <= matchd386d;
	-- d388d
	sted388d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord388d,
			Enable=>Enabled388d,
			match=>matchd388d,
			run=>run);

	Enabled388d <= matchd387d;
	-- d389d
	sted389d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord389d,
			Enable=>Enabled389d,
			match=>matchd389d,
			run=>run);

	Enabled389d <= matchd388d;
	-- d390d
	sted390d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord390d,
			Enable=>Enabled390d,
			match=>matchd390d,
			run=>run);

	Enabled390d <= matchd389d;
	-- d391d
	sted391d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord391d,
			Enable=>Enabled391d,
			match=>matchd391d,
			run=>run);

	-- d392d
	sted392d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord392d,
			Enable=>Enabled392d,
			match=>matchd392d,
			run=>run);

	Enabled392d <= matchd392d OR matchd391d;
	-- d393d
	sted393d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord393d,
			Enable=>Enabled393d,
			match=>matchd393d,
			run=>run);

	Enabled393d <= matchd392d;
	-- d394d
	sted394d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord394d,
			Enable=>Enabled394d,
			match=>matchd394d,
			run=>run);

	Enabled394d <= matchd394d OR matchd393d;
	-- d395d
	sted395d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord395d,
			Enable=>Enabled395d,
			match=>matchd395d,
			run=>run);

	Enabled395d <= matchd394d;
	-- d396d
	sted396d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord396d,
			Enable=>Enabled396d,
			match=>matchd396d,
			run=>run);

	Enabled396d <= matchd396d OR matchd395d;
	-- d397d
	sted397d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord397d,
			Enable=>Enabled397d,
			match=>matchd397d,
			run=>run);

	Enabled397d <= matchd396d;
	-- d398d
	sted398d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord398d,
			Enable=>Enabled398d,
			match=>matchd398d,
			run=>run);

	Enabled398d <= matchd397d;
	-- d399d
	sted399d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord399d,
			Enable=>Enabled399d,
			match=>matchd399d,
			run=>run);

	Enabled399d <= matchd398d;
	-- d400d
	sted400d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord400d,
			Enable=>Enabled400d,
			match=>matchd400d,
			run=>run);

	Enabled400d <= matchd399d;
	-- d401d
	sted401d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord401d,
			Enable=>Enabled401d,
			match=>matchd401d,
			run=>run);

	Enabled401d <= matchd400d;
	-- d402d
	sted402d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord402d,
			Enable=>Enabled402d,
			match=>matchd402d,
			run=>run);

	Enabled402d <= matchd401d OR matchd402d;
	-- d403d
	sted403d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord403d,
			Enable=>Enabled403d,
			match=>matchd403d,
			run=>run);

	Enabled403d <= matchd402d;
	-- d404d
	sted404d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord404d,
			Enable=>Enabled404d,
			match=>matchd404d,
			run=>run);

	Enabled404d <= matchd403d OR matchd404d;
	-- d405d
	sted405d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord405d,
			Enable=>Enabled405d,
			match=>matchd405d,
			run=>run);

	Enabled405d <= matchd404d;
	-- d406d
	sted406d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord406d,
			Enable=>Enabled406d,
			match=>matchd406d,
			run=>run);

	Enabled406d <= matchd405d OR matchd406d;
	-- d407d
	sted407d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord407d,
			Enable=>Enabled407d,
			match=>matchd407d,
			run=>run);

	Enabled407d <= matchd406d;
	-- d408d
	sted408d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord408d,
			Enable=>Enabled408d,
			match=>matchd408d,
			run=>run);

	Enabled408d <= matchd407d;
	-- d409d
	sted409d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord409d,
			Enable=>Enabled409d,
			match=>matchd409d,
			run=>run);

	Enabled409d <= matchd408d;
	-- d410d
	sted410d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord410d,
			Enable=>Enabled410d,
			match=>matchd410d,
			run=>run);

	Enabled410d <= matchd409d;
	-- d411d
	sted411d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord411d,
			Enable=>Enabled411d,
			match=>matchd411d,
			run=>run);

	Enabled411d <= matchd410d;
	-- d412d
	sted412d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord412d,
			Enable=>Enabled412d,
			match=>matchd412d,
			run=>run);

	-- d413d
	sted413d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord413d,
			Enable=>Enabled413d,
			match=>matchd413d,
			run=>run);

	Enabled413d <= matchd413d OR matchd412d;
	-- d414d
	sted414d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord414d,
			Enable=>Enabled414d,
			match=>matchd414d,
			run=>run);

	Enabled414d <= matchd413d;
	-- d415d
	sted415d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord415d,
			Enable=>Enabled415d,
			match=>matchd415d,
			run=>run);

	Enabled415d <= matchd414d OR matchd415d;
	-- d416d
	sted416d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord416d,
			Enable=>Enabled416d,
			match=>matchd416d,
			run=>run);

	Enabled416d <= matchd415d;
	-- d417d
	sted417d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord417d,
			Enable=>Enabled417d,
			match=>matchd417d,
			run=>run);

	Enabled417d <= matchd417d OR matchd416d;
	-- d418d
	sted418d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord418d,
			Enable=>Enabled418d,
			match=>matchd418d,
			run=>run);

	Enabled418d <= matchd417d;
	-- d419d
	sted419d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord419d,
			Enable=>Enabled419d,
			match=>matchd419d,
			run=>run);

	Enabled419d <= matchd419d OR matchd418d;
	-- d420d
	sted420d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord420d,
			Enable=>Enabled420d,
			match=>matchd420d,
			run=>run);

	Enabled420d <= matchd419d;
	-- d421d
	sted421d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord421d,
			Enable=>Enabled421d,
			match=>matchd421d,
			run=>run);

	Enabled421d <= matchd420d OR matchd421d;
	-- d422d
	sted422d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord422d,
			Enable=>Enabled422d,
			match=>matchd422d,
			run=>run);

	Enabled422d <= matchd421d;
	-- d423d
	sted423d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord423d,
			Enable=>Enabled423d,
			match=>matchd423d,
			run=>run);

	Enabled423d <= matchd422d;
	-- d424d
	sted424d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord424d,
			Enable=>Enabled424d,
			match=>matchd424d,
			run=>run);

	Enabled424d <= matchd423d;
	-- d425d
	sted425d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord425d,
			Enable=>Enabled425d,
			match=>matchd425d,
			run=>run);

	Enabled425d <= matchd424d;
	-- d426d
	sted426d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord426d,
			Enable=>Enabled426d,
			match=>matchd426d,
			run=>run);

	Enabled426d <= matchd425d;
	-- d427d
	sted427d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord427d,
			Enable=>Enabled427d,
			match=>matchd427d,
			run=>run);

	Enabled427d <= matchd427d OR matchd426d;
	-- d428d
	sted428d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord428d,
			Enable=>Enabled428d,
			match=>matchd428d,
			run=>run);

	Enabled428d <= matchd427d;
	-- d429d
	sted429d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord429d,
			Enable=>Enabled429d,
			match=>matchd429d,
			run=>run);

	Enabled429d <= matchd428d;
	-- d430d
	sted430d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord430d,
			Enable=>Enabled430d,
			match=>matchd430d,
			run=>run);

	Enabled430d <= matchd429d;
	-- d431d
	sted431d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord431d,
			Enable=>Enabled431d,
			match=>matchd431d,
			run=>run);

	Enabled431d <= matchd430d;
	-- d432d
	sted432d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord432d,
			Enable=>Enabled432d,
			match=>matchd432d,
			run=>run);

	Enabled432d <= matchd431d;
	-- d434d
	sted434d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord434d,
			Enable=>Enabled434d,
			match=>matchd434d,
			run=>run);

	-- d435d
	sted435d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord435d,
			Enable=>Enabled435d,
			match=>matchd435d,
			run=>run);

	Enabled435d <= matchd435d OR matchd434d;
	-- d436d
	sted436d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord436d,
			Enable=>Enabled436d,
			match=>matchd436d,
			run=>run);

	Enabled436d <= matchd435d;
	-- d437d
	sted437d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord437d,
			Enable=>Enabled437d,
			match=>matchd437d,
			run=>run);

	Enabled437d <= matchd436d;
	-- d438d
	sted438d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord438d,
			Enable=>Enabled438d,
			match=>matchd438d,
			run=>run);

	Enabled438d <= matchd437d;
	-- d439d
	sted439d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord439d,
			Enable=>Enabled439d,
			match=>matchd439d,
			run=>run);

	Enabled439d <= matchd438d;
	-- d440d
	sted440d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord440d,
			Enable=>Enabled440d,
			match=>matchd440d,
			run=>run);

	Enabled440d <= matchd439d OR matchd440d;
	-- d441d
	sted441d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord441d,
			Enable=>Enabled441d,
			match=>matchd441d,
			run=>run);

	Enabled441d <= matchd440d;
	-- d442d
	sted442d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord442d,
			Enable=>Enabled442d,
			match=>matchd442d,
			run=>run);

	Enabled442d <= matchd441d;
	-- d443d
	sted443d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord443d,
			Enable=>Enabled443d,
			match=>matchd443d,
			run=>run);

	Enabled443d <= matchd442d;
	-- d444d
	sted444d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord444d,
			Enable=>Enabled444d,
			match=>matchd444d,
			run=>run);

	reports(21) <= matchd444d;
	Enabled444d <= matchd443d;
	-- d445d
	sted445d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord445d,
			Enable=>Enabled445d,
			match=>matchd445d,
			run=>run);

	-- d446d
	sted446d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord446d,
			Enable=>Enabled446d,
			match=>matchd446d,
			run=>run);

	Enabled446d <= matchd445d OR matchd446d;
	-- d447d
	sted447d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord447d,
			Enable=>Enabled447d,
			match=>matchd447d,
			run=>run);

	Enabled447d <= matchd446d;
	-- d448d
	sted448d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord448d,
			Enable=>Enabled448d,
			match=>matchd448d,
			run=>run);

	Enabled448d <= matchd447d;
	-- d449d
	sted449d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord449d,
			Enable=>Enabled449d,
			match=>matchd449d,
			run=>run);

	Enabled449d <= matchd448d;
	-- d450d
	sted450d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord450d,
			Enable=>Enabled450d,
			match=>matchd450d,
			run=>run);

	Enabled450d <= matchd449d;
	-- d451d
	sted451d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord451d,
			Enable=>Enabled451d,
			match=>matchd451d,
			run=>run);

	Enabled451d <= matchd450d OR matchd451d;
	-- d452d
	sted452d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord452d,
			Enable=>Enabled452d,
			match=>matchd452d,
			run=>run);

	Enabled452d <= matchd451d;
	-- d453d
	sted453d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord453d,
			Enable=>Enabled453d,
			match=>matchd453d,
			run=>run);

	Enabled453d <= matchd453d OR matchd452d;
	-- d454d
	sted454d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord454d,
			Enable=>Enabled454d,
			match=>matchd454d,
			run=>run);

	Enabled454d <= matchd453d;
	-- d455d
	sted455d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord455d,
			Enable=>Enabled455d,
			match=>matchd455d,
			run=>run);

	Enabled455d <= matchd455d OR matchd454d;
	-- d456d
	sted456d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord456d,
			Enable=>Enabled456d,
			match=>matchd456d,
			run=>run);

	Enabled456d <= matchd455d;
	-- d457d
	sted457d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord457d,
			Enable=>Enabled457d,
			match=>matchd457d,
			run=>run);

	Enabled457d <= matchd457d OR matchd456d;
	-- d458d
	sted458d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord458d,
			Enable=>Enabled458d,
			match=>matchd458d,
			run=>run);

	Enabled458d <= matchd457d;
	-- d459d
	sted459d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord459d,
			Enable=>Enabled459d,
			match=>matchd459d,
			run=>run);

	Enabled459d <= matchd459d OR matchd458d;
	-- d460d
	sted460d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord460d,
			Enable=>Enabled460d,
			match=>matchd460d,
			run=>run);

	Enabled460d <= matchd459d;
	-- d461d
	sted461d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord461d,
			Enable=>Enabled461d,
			match=>matchd461d,
			run=>run);

	Enabled461d <= matchd460d;
	-- d462d
	sted462d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord462d,
			Enable=>Enabled462d,
			match=>matchd462d,
			run=>run);

	Enabled462d <= matchd461d;
	-- d463d
	sted463d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord463d,
			Enable=>Enabled463d,
			match=>matchd463d,
			run=>run);

	Enabled463d <= matchd462d;
	-- d464d
	sted464d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord464d,
			Enable=>Enabled464d,
			match=>matchd464d,
			run=>run);

	Enabled464d <= matchd463d;
	-- d465d
	sted465d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord465d,
			Enable=>Enabled465d,
			match=>matchd465d,
			run=>run);

	-- d466d
	sted466d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord466d,
			Enable=>Enabled466d,
			match=>matchd466d,
			run=>run);

	Enabled466d <= matchd466d OR matchd465d;
	-- d467d
	sted467d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord467d,
			Enable=>Enabled467d,
			match=>matchd467d,
			run=>run);

	Enabled467d <= matchd466d;
	-- d468d
	sted468d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord468d,
			Enable=>Enabled468d,
			match=>matchd468d,
			run=>run);

	Enabled468d <= matchd467d OR matchd468d;
	-- d469d
	sted469d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord469d,
			Enable=>Enabled469d,
			match=>matchd469d,
			run=>run);

	Enabled469d <= matchd468d;
	-- d470d
	sted470d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord470d,
			Enable=>Enabled470d,
			match=>matchd470d,
			run=>run);

	Enabled470d <= matchd470d OR matchd469d;
	-- d471d
	sted471d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord471d,
			Enable=>Enabled471d,
			match=>matchd471d,
			run=>run);

	Enabled471d <= matchd470d;
	-- d472d
	sted472d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord472d,
			Enable=>Enabled472d,
			match=>matchd472d,
			run=>run);

	Enabled472d <= matchd471d;
	-- d473d
	sted473d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord473d,
			Enable=>Enabled473d,
			match=>matchd473d,
			run=>run);

	Enabled473d <= matchd472d;
	-- d474d
	sted474d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord474d,
			Enable=>Enabled474d,
			match=>matchd474d,
			run=>run);

	Enabled474d <= matchd473d;
	-- d475d
	sted475d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord475d,
			Enable=>Enabled475d,
			match=>matchd475d,
			run=>run);

	Enabled475d <= matchd475d OR matchd474d;
	-- d476d
	sted476d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord476d,
			Enable=>Enabled476d,
			match=>matchd476d,
			run=>run);

	Enabled476d <= matchd475d;
	-- d477d
	sted477d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord477d,
			Enable=>Enabled477d,
			match=>matchd477d,
			run=>run);

	Enabled477d <= matchd477d OR matchd476d;
	-- d478d
	sted478d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord478d,
			Enable=>Enabled478d,
			match=>matchd478d,
			run=>run);

	Enabled478d <= matchd477d;
	-- d479d
	sted479d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord479d,
			Enable=>Enabled479d,
			match=>matchd479d,
			run=>run);

	Enabled479d <= matchd479d OR matchd478d;
	-- d480d
	sted480d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord480d,
			Enable=>Enabled480d,
			match=>matchd480d,
			run=>run);

	Enabled480d <= matchd479d;
	-- d481d
	sted481d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord481d,
			Enable=>Enabled481d,
			match=>matchd481d,
			run=>run);

	Enabled481d <= matchd480d;
	-- d482d
	sted482d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord482d,
			Enable=>Enabled482d,
			match=>matchd482d,
			run=>run);

	Enabled482d <= matchd481d;
	-- d483d
	sted483d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord483d,
			Enable=>Enabled483d,
			match=>matchd483d,
			run=>run);

	Enabled483d <= matchd482d;
	-- d484d
	sted484d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord484d,
			Enable=>Enabled484d,
			match=>matchd484d,
			run=>run);

	Enabled484d <= matchd483d;
	-- d485d
	sted485d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord485d,
			Enable=>Enabled485d,
			match=>matchd485d,
			run=>run);

	-- d486d
	sted486d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord486d,
			Enable=>Enabled486d,
			match=>matchd486d,
			run=>run);

	Enabled486d <= matchd485d OR matchd486d;
	-- d487d
	sted487d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord487d,
			Enable=>Enabled487d,
			match=>matchd487d,
			run=>run);

	Enabled487d <= matchd486d;
	-- d488d
	sted488d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord488d,
			Enable=>Enabled488d,
			match=>matchd488d,
			run=>run);

	Enabled488d <= matchd487d OR matchd488d;
	-- d489d
	sted489d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord489d,
			Enable=>Enabled489d,
			match=>matchd489d,
			run=>run);

	Enabled489d <= matchd488d;
	-- d490d
	sted490d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord490d,
			Enable=>Enabled490d,
			match=>matchd490d,
			run=>run);

	Enabled490d <= matchd489d OR matchd490d;
	-- d491d
	sted491d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord491d,
			Enable=>Enabled491d,
			match=>matchd491d,
			run=>run);

	Enabled491d <= matchd490d;
	-- d492d
	sted492d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord492d,
			Enable=>Enabled492d,
			match=>matchd492d,
			run=>run);

	Enabled492d <= matchd492d OR matchd491d;
	-- d493d
	sted493d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord493d,
			Enable=>Enabled493d,
			match=>matchd493d,
			run=>run);

	Enabled493d <= matchd492d;
	-- d494d
	sted494d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord494d,
			Enable=>Enabled494d,
			match=>matchd494d,
			run=>run);

	Enabled494d <= matchd494d OR matchd493d;
	-- d495d
	sted495d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord495d,
			Enable=>Enabled495d,
			match=>matchd495d,
			run=>run);

	Enabled495d <= matchd494d;
	-- d496d
	sted496d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord496d,
			Enable=>Enabled496d,
			match=>matchd496d,
			run=>run);

	Enabled496d <= matchd495d;
	-- d497d
	sted497d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord497d,
			Enable=>Enabled497d,
			match=>matchd497d,
			run=>run);

	Enabled497d <= matchd496d;
	-- d498d
	sted498d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord498d,
			Enable=>Enabled498d,
			match=>matchd498d,
			run=>run);

	Enabled498d <= matchd497d;
	-- d499d
	sted499d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord499d,
			Enable=>Enabled499d,
			match=>matchd499d,
			run=>run);

	Enabled499d <= matchd499d OR matchd498d;
	-- d500d
	sted500d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord500d,
			Enable=>Enabled500d,
			match=>matchd500d,
			run=>run);

	Enabled500d <= matchd499d;
	-- d501d
	sted501d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord501d,
			Enable=>Enabled501d,
			match=>matchd501d,
			run=>run);

	Enabled501d <= matchd500d;
	-- d502d
	sted502d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord502d,
			Enable=>Enabled502d,
			match=>matchd502d,
			run=>run);

	Enabled502d <= matchd501d;
	-- d503d
	sted503d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord503d,
			Enable=>Enabled503d,
			match=>matchd503d,
			run=>run);

	Enabled503d <= matchd502d;
	-- d504d
	sted504d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord504d,
			Enable=>Enabled504d,
			match=>matchd504d,
			run=>run);

	Enabled504d <= matchd503d;
	-- d506d
	sted506d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord506d,
			Enable=>Enabled506d,
			match=>matchd506d,
			run=>run);

	-- d507d
	sted507d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord507d,
			Enable=>Enabled507d,
			match=>matchd507d,
			run=>run);

	Enabled507d <= matchd506d;
	-- d508d
	sted508d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord508d,
			Enable=>Enabled508d,
			match=>matchd508d,
			run=>run);

	Enabled508d <= matchd507d;
	-- d509d
	sted509d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord509d,
			Enable=>Enabled509d,
			match=>matchd509d,
			run=>run);

	Enabled509d <= matchd508d;
	-- d510d
	sted510d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord510d,
			Enable=>Enabled510d,
			match=>matchd510d,
			run=>run);

	Enabled510d <= matchd509d;
	-- d511d
	sted511d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord511d,
			Enable=>Enabled511d,
			match=>matchd511d,
			run=>run);

	Enabled511d <= matchd510d;
	-- d512d
	sted512d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord512d,
			Enable=>Enabled512d,
			match=>matchd512d,
			run=>run);

	Enabled512d <= matchd511d;
	-- d513d
	sted513d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord513d,
			Enable=>Enabled513d,
			match=>matchd513d,
			run=>run);

	Enabled513d <= matchd512d OR matchd513d;
	-- d514d
	sted514d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord514d,
			Enable=>Enabled514d,
			match=>matchd514d,
			run=>run);

	Enabled514d <= matchd513d;
	-- d515d
	sted515d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord515d,
			Enable=>Enabled515d,
			match=>matchd515d,
			run=>run);

	Enabled515d <= matchd514d OR matchd515d;
	-- d516d
	sted516d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord516d,
			Enable=>Enabled516d,
			match=>matchd516d,
			run=>run);

	Enabled516d <= matchd515d;
	-- d517d
	sted517d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord517d,
			Enable=>Enabled517d,
			match=>matchd517d,
			run=>run);

	Enabled517d <= matchd516d;
	-- d518d
	sted518d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord518d,
			Enable=>Enabled518d,
			match=>matchd518d,
			run=>run);

	Enabled518d <= matchd517d;
	-- d519d
	sted519d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord519d,
			Enable=>Enabled519d,
			match=>matchd519d,
			run=>run);

	Enabled519d <= matchd518d;
	-- d520d
	sted520d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord520d,
			Enable=>Enabled520d,
			match=>matchd520d,
			run=>run);

	Enabled520d <= matchd519d OR matchd520d;
	-- d521d
	sted521d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord521d,
			Enable=>Enabled521d,
			match=>matchd521d,
			run=>run);

	reports(22) <= matchd521d;
	Enabled521d <= matchd520d;
	-- d522d
	sted522d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord522d,
			Enable=>Enabled522d,
			match=>matchd522d,
			run=>run);

	-- d523d
	sted523d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord523d,
			Enable=>Enabled523d,
			match=>matchd523d,
			run=>run);

	Enabled523d <= matchd523d OR matchd522d;
	-- d524d
	sted524d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord524d,
			Enable=>Enabled524d,
			match=>matchd524d,
			run=>run);

	Enabled524d <= matchd523d;
	-- d525d
	sted525d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord525d,
			Enable=>Enabled525d,
			match=>matchd525d,
			run=>run);

	Enabled525d <= matchd524d OR matchd525d;
	-- d526d
	sted526d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord526d,
			Enable=>Enabled526d,
			match=>matchd526d,
			run=>run);

	Enabled526d <= matchd525d;
	-- d527d
	sted527d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord527d,
			Enable=>Enabled527d,
			match=>matchd527d,
			run=>run);

	Enabled527d <= matchd526d OR matchd527d;
	-- d528d
	sted528d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord528d,
			Enable=>Enabled528d,
			match=>matchd528d,
			run=>run);

	Enabled528d <= matchd527d;
	-- d529d
	sted529d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord529d,
			Enable=>Enabled529d,
			match=>matchd529d,
			run=>run);

	Enabled529d <= matchd528d;
	-- d530d
	sted530d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord530d,
			Enable=>Enabled530d,
			match=>matchd530d,
			run=>run);

	Enabled530d <= matchd529d;
	-- d531d
	sted531d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord531d,
			Enable=>Enabled531d,
			match=>matchd531d,
			run=>run);

	Enabled531d <= matchd530d;
	-- d532d
	sted532d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord532d,
			Enable=>Enabled532d,
			match=>matchd532d,
			run=>run);

	Enabled532d <= matchd531d OR matchd532d;
	-- d533d
	sted533d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord533d,
			Enable=>Enabled533d,
			match=>matchd533d,
			run=>run);

	Enabled533d <= matchd532d;
	-- d534d
	sted534d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord534d,
			Enable=>Enabled534d,
			match=>matchd534d,
			run=>run);

	Enabled534d <= matchd533d;
	-- d535d
	sted535d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord535d,
			Enable=>Enabled535d,
			match=>matchd535d,
			run=>run);

	Enabled535d <= matchd534d;
	-- d536d
	sted536d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord536d,
			Enable=>Enabled536d,
			match=>matchd536d,
			run=>run);

	Enabled536d <= matchd535d;
	-- d537d
	sted537d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord537d,
			Enable=>Enabled537d,
			match=>matchd537d,
			run=>run);

	Enabled537d <= matchd536d;
	-- d538d
	sted538d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord538d,
			Enable=>Enabled538d,
			match=>matchd538d,
			run=>run);

	-- d539d
	sted539d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord539d,
			Enable=>Enabled539d,
			match=>matchd539d,
			run=>run);

	Enabled539d <= matchd538d OR matchd539d;
	-- d540d
	sted540d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord540d,
			Enable=>Enabled540d,
			match=>matchd540d,
			run=>run);

	Enabled540d <= matchd539d;
	-- d541d
	sted541d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord541d,
			Enable=>Enabled541d,
			match=>matchd541d,
			run=>run);

	Enabled541d <= matchd540d;
	-- d542d
	sted542d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord542d,
			Enable=>Enabled542d,
			match=>matchd542d,
			run=>run);

	Enabled542d <= matchd541d;
	-- d543d
	sted543d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord543d,
			Enable=>Enabled543d,
			match=>matchd543d,
			run=>run);

	Enabled543d <= matchd542d;
	-- d544d
	sted544d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord544d,
			Enable=>Enabled544d,
			match=>matchd544d,
			run=>run);

	Enabled544d <= matchd543d OR matchd544d;
	-- d545d
	sted545d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord545d,
			Enable=>Enabled545d,
			match=>matchd545d,
			run=>run);

	Enabled545d <= matchd544d;
	-- d546d
	sted546d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord546d,
			Enable=>Enabled546d,
			match=>matchd546d,
			run=>run);

	Enabled546d <= matchd546d OR matchd545d;
	-- d547d
	sted547d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord547d,
			Enable=>Enabled547d,
			match=>matchd547d,
			run=>run);

	Enabled547d <= matchd546d;
	-- d548d
	sted548d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord548d,
			Enable=>Enabled548d,
			match=>matchd548d,
			run=>run);

	Enabled548d <= matchd548d OR matchd547d;
	-- d549d
	sted549d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord549d,
			Enable=>Enabled549d,
			match=>matchd549d,
			run=>run);

	Enabled549d <= matchd548d;
	-- d550d
	sted550d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord550d,
			Enable=>Enabled550d,
			match=>matchd550d,
			run=>run);

	Enabled550d <= matchd549d;
	-- d551d
	sted551d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord551d,
			Enable=>Enabled551d,
			match=>matchd551d,
			run=>run);

	Enabled551d <= matchd550d;
	-- d552d
	sted552d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord552d,
			Enable=>Enabled552d,
			match=>matchd552d,
			run=>run);

	Enabled552d <= matchd551d;
	-- d553d
	sted553d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord553d,
			Enable=>Enabled553d,
			match=>matchd553d,
			run=>run);

	Enabled553d <= matchd552d;
	-- d555d
	sted555d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord555d,
			Enable=>Enabled555d,
			match=>matchd555d,
			run=>run);

	-- d556d
	sted556d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord556d,
			Enable=>Enabled556d,
			match=>matchd556d,
			run=>run);

	Enabled556d <= matchd556d OR matchd555d;
	-- d557d
	sted557d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord557d,
			Enable=>Enabled557d,
			match=>matchd557d,
			run=>run);

	Enabled557d <= matchd556d;
	-- d558d
	sted558d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord558d,
			Enable=>Enabled558d,
			match=>matchd558d,
			run=>run);

	Enabled558d <= matchd557d;
	-- d559d
	sted559d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord559d,
			Enable=>Enabled559d,
			match=>matchd559d,
			run=>run);

	Enabled559d <= matchd558d;
	-- d560d
	sted560d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord560d,
			Enable=>Enabled560d,
			match=>matchd560d,
			run=>run);

	Enabled560d <= matchd559d;
	-- d561d
	sted561d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord561d,
			Enable=>Enabled561d,
			match=>matchd561d,
			run=>run);

	Enabled561d <= matchd561d OR matchd560d;
	-- d562d
	sted562d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord562d,
			Enable=>Enabled562d,
			match=>matchd562d,
			run=>run);

	Enabled562d <= matchd561d;
	-- d563d
	sted563d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord563d,
			Enable=>Enabled563d,
			match=>matchd563d,
			run=>run);

	Enabled563d <= matchd562d;
	-- d564d
	sted564d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord564d,
			Enable=>Enabled564d,
			match=>matchd564d,
			run=>run);

	Enabled564d <= matchd563d;
	-- d565d
	sted565d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord565d,
			Enable=>Enabled565d,
			match=>matchd565d,
			run=>run);

	reports(23) <= matchd565d;
	Enabled565d <= matchd564d;
	-- d566d
	sted566d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord566d,
			Enable=>Enabled566d,
			match=>matchd566d,
			run=>run);

	-- d567d
	sted567d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord567d,
			Enable=>Enabled567d,
			match=>matchd567d,
			run=>run);

	Enabled567d <= matchd567d OR matchd566d;
	-- d568d
	sted568d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord568d,
			Enable=>Enabled568d,
			match=>matchd568d,
			run=>run);

	Enabled568d <= matchd567d;
	-- d569d
	sted569d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord569d,
			Enable=>Enabled569d,
			match=>matchd569d,
			run=>run);

	Enabled569d <= matchd568d;
	-- d570d
	sted570d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord570d,
			Enable=>Enabled570d,
			match=>matchd570d,
			run=>run);

	Enabled570d <= matchd569d;
	-- d571d
	sted571d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord571d,
			Enable=>Enabled571d,
			match=>matchd571d,
			run=>run);

	Enabled571d <= matchd570d;
	-- d572d
	sted572d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord572d,
			Enable=>Enabled572d,
			match=>matchd572d,
			run=>run);

	Enabled572d <= matchd571d OR matchd572d;
	-- d573d
	sted573d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord573d,
			Enable=>Enabled573d,
			match=>matchd573d,
			run=>run);

	Enabled573d <= matchd572d;
	-- d574d
	sted574d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord574d,
			Enable=>Enabled574d,
			match=>matchd574d,
			run=>run);

	Enabled574d <= matchd573d OR matchd574d;
	-- d575d
	sted575d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord575d,
			Enable=>Enabled575d,
			match=>matchd575d,
			run=>run);

	Enabled575d <= matchd574d;
	-- d576d
	sted576d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord576d,
			Enable=>Enabled576d,
			match=>matchd576d,
			run=>run);

	Enabled576d <= matchd575d OR matchd576d;
	-- d577d
	sted577d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord577d,
			Enable=>Enabled577d,
			match=>matchd577d,
			run=>run);

	Enabled577d <= matchd576d;
	-- d578d
	sted578d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord578d,
			Enable=>Enabled578d,
			match=>matchd578d,
			run=>run);

	Enabled578d <= matchd577d OR matchd578d;
	-- d579d
	sted579d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord579d,
			Enable=>Enabled579d,
			match=>matchd579d,
			run=>run);

	Enabled579d <= matchd578d;
	-- d580d
	sted580d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord580d,
			Enable=>Enabled580d,
			match=>matchd580d,
			run=>run);

	Enabled580d <= matchd580d OR matchd579d;
	-- d581d
	sted581d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord581d,
			Enable=>Enabled581d,
			match=>matchd581d,
			run=>run);

	Enabled581d <= matchd580d;
	-- d582d
	sted582d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord582d,
			Enable=>Enabled582d,
			match=>matchd582d,
			run=>run);

	Enabled582d <= matchd581d;
	-- d583d
	sted583d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord583d,
			Enable=>Enabled583d,
			match=>matchd583d,
			run=>run);

	Enabled583d <= matchd582d;
	-- d584d
	sted584d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord584d,
			Enable=>Enabled584d,
			match=>matchd584d,
			run=>run);

	Enabled584d <= matchd583d;
	-- d585d
	sted585d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord585d,
			Enable=>Enabled585d,
			match=>matchd585d,
			run=>run);

	Enabled585d <= matchd584d;
	-- d586d
	sted586d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord586d,
			Enable=>Enabled586d,
			match=>matchd586d,
			run=>run);

	-- d587d
	sted587d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord587d,
			Enable=>Enabled587d,
			match=>matchd587d,
			run=>run);

	Enabled587d <= matchd587d OR matchd586d;
	-- d588d
	sted588d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord588d,
			Enable=>Enabled588d,
			match=>matchd588d,
			run=>run);

	Enabled588d <= matchd587d;
	-- d589d
	sted589d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord589d,
			Enable=>Enabled589d,
			match=>matchd589d,
			run=>run);

	Enabled589d <= matchd589d OR matchd588d;
	-- d590d
	sted590d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord590d,
			Enable=>Enabled590d,
			match=>matchd590d,
			run=>run);

	Enabled590d <= matchd589d;
	-- d591d
	sted591d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord591d,
			Enable=>Enabled591d,
			match=>matchd591d,
			run=>run);

	Enabled591d <= matchd590d OR matchd591d;
	-- d592d
	sted592d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord592d,
			Enable=>Enabled592d,
			match=>matchd592d,
			run=>run);

	Enabled592d <= matchd591d;
	-- d593d
	sted593d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord593d,
			Enable=>Enabled593d,
			match=>matchd593d,
			run=>run);

	Enabled593d <= matchd592d;
	-- d594d
	sted594d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord594d,
			Enable=>Enabled594d,
			match=>matchd594d,
			run=>run);

	Enabled594d <= matchd593d;
	-- d595d
	sted595d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord595d,
			Enable=>Enabled595d,
			match=>matchd595d,
			run=>run);

	Enabled595d <= matchd594d;
	-- d596d
	sted596d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord596d,
			Enable=>Enabled596d,
			match=>matchd596d,
			run=>run);

	Enabled596d <= matchd595d OR matchd596d;
	-- d597d
	sted597d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord597d,
			Enable=>Enabled597d,
			match=>matchd597d,
			run=>run);

	Enabled597d <= matchd596d;
	-- d598d
	sted598d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord598d,
			Enable=>Enabled598d,
			match=>matchd598d,
			run=>run);

	Enabled598d <= matchd598d OR matchd597d;
	-- d599d
	sted599d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord599d,
			Enable=>Enabled599d,
			match=>matchd599d,
			run=>run);

	Enabled599d <= matchd598d;
	-- d600d
	sted600d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord600d,
			Enable=>Enabled600d,
			match=>matchd600d,
			run=>run);

	Enabled600d <= matchd599d OR matchd600d;
	-- d601d
	sted601d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord601d,
			Enable=>Enabled601d,
			match=>matchd601d,
			run=>run);

	Enabled601d <= matchd600d;
	-- d602d
	sted602d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord602d,
			Enable=>Enabled602d,
			match=>matchd602d,
			run=>run);

	Enabled602d <= matchd601d;
	-- d603d
	sted603d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord603d,
			Enable=>Enabled603d,
			match=>matchd603d,
			run=>run);

	Enabled603d <= matchd602d;
	-- d604d
	sted604d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord604d,
			Enable=>Enabled604d,
			match=>matchd604d,
			run=>run);

	Enabled604d <= matchd603d;
	-- d605d
	sted605d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord605d,
			Enable=>Enabled605d,
			match=>matchd605d,
			run=>run);

	Enabled605d <= matchd604d;
	-- d606d
	sted606d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord606d,
			Enable=>Enabled606d,
			match=>matchd606d,
			run=>run);

	-- d607d
	sted607d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord607d,
			Enable=>Enabled607d,
			match=>matchd607d,
			run=>run);

	Enabled607d <= matchd606d OR matchd607d;
	-- d608d
	sted608d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord608d,
			Enable=>Enabled608d,
			match=>matchd608d,
			run=>run);

	Enabled608d <= matchd607d;
	-- d609d
	sted609d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord609d,
			Enable=>Enabled609d,
			match=>matchd609d,
			run=>run);

	Enabled609d <= matchd608d OR matchd609d;
	-- d610d
	sted610d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord610d,
			Enable=>Enabled610d,
			match=>matchd610d,
			run=>run);

	Enabled610d <= matchd609d;
	-- d611d
	sted611d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord611d,
			Enable=>Enabled611d,
			match=>matchd611d,
			run=>run);

	Enabled611d <= matchd611d OR matchd610d;
	-- d612d
	sted612d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord612d,
			Enable=>Enabled612d,
			match=>matchd612d,
			run=>run);

	Enabled612d <= matchd611d;
	-- d613d
	sted613d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord613d,
			Enable=>Enabled613d,
			match=>matchd613d,
			run=>run);

	Enabled613d <= matchd612d OR matchd613d;
	-- d614d
	sted614d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord614d,
			Enable=>Enabled614d,
			match=>matchd614d,
			run=>run);

	Enabled614d <= matchd613d;
	-- d615d
	sted615d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord615d,
			Enable=>Enabled615d,
			match=>matchd615d,
			run=>run);

	Enabled615d <= matchd614d OR matchd615d;
	-- d616d
	sted616d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord616d,
			Enable=>Enabled616d,
			match=>matchd616d,
			run=>run);

	Enabled616d <= matchd615d;
	-- d617d
	sted617d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord617d,
			Enable=>Enabled617d,
			match=>matchd617d,
			run=>run);

	Enabled617d <= matchd616d;
	-- d618d
	sted618d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord618d,
			Enable=>Enabled618d,
			match=>matchd618d,
			run=>run);

	Enabled618d <= matchd617d;
	-- d619d
	sted619d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord619d,
			Enable=>Enabled619d,
			match=>matchd619d,
			run=>run);

	Enabled619d <= matchd618d;
	-- d620d
	sted620d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord620d,
			Enable=>Enabled620d,
			match=>matchd620d,
			run=>run);

	Enabled620d <= matchd619d OR matchd620d;
	-- d621d
	sted621d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord621d,
			Enable=>Enabled621d,
			match=>matchd621d,
			run=>run);

	Enabled621d <= matchd620d;
	-- d622d
	sted622d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord622d,
			Enable=>Enabled622d,
			match=>matchd622d,
			run=>run);

	Enabled622d <= matchd621d;
	-- d623d
	sted623d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord623d,
			Enable=>Enabled623d,
			match=>matchd623d,
			run=>run);

	Enabled623d <= matchd622d;
	-- d624d
	sted624d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord624d,
			Enable=>Enabled624d,
			match=>matchd624d,
			run=>run);

	Enabled624d <= matchd623d;
	-- d625d
	sted625d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord625d,
			Enable=>Enabled625d,
			match=>matchd625d,
			run=>run);

	Enabled625d <= matchd624d;
	-- d627d
	sted627d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord627d,
			Enable=>Enabled627d,
			match=>matchd627d,
			run=>run);

	-- d628d
	sted628d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord628d,
			Enable=>Enabled628d,
			match=>matchd628d,
			run=>run);

	Enabled628d <= matchd628d OR matchd627d;
	-- d629d
	sted629d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord629d,
			Enable=>Enabled629d,
			match=>matchd629d,
			run=>run);

	Enabled629d <= matchd628d;
	-- d630d
	sted630d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord630d,
			Enable=>Enabled630d,
			match=>matchd630d,
			run=>run);

	Enabled630d <= matchd629d;
	-- d631d
	sted631d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord631d,
			Enable=>Enabled631d,
			match=>matchd631d,
			run=>run);

	Enabled631d <= matchd630d;
	-- d632d
	sted632d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord632d,
			Enable=>Enabled632d,
			match=>matchd632d,
			run=>run);

	Enabled632d <= matchd631d;
	-- d633d
	sted633d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord633d,
			Enable=>Enabled633d,
			match=>matchd633d,
			run=>run);

	Enabled633d <= matchd632d;
	-- d634d
	sted634d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord634d,
			Enable=>Enabled634d,
			match=>matchd634d,
			run=>run);

	Enabled634d <= matchd634d OR matchd633d;
	-- d635d
	sted635d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord635d,
			Enable=>Enabled635d,
			match=>matchd635d,
			run=>run);

	Enabled635d <= matchd634d;
	-- d636d
	sted636d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord636d,
			Enable=>Enabled636d,
			match=>matchd636d,
			run=>run);

	Enabled636d <= matchd635d;
	-- d637d
	sted637d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord637d,
			Enable=>Enabled637d,
			match=>matchd637d,
			run=>run);

	Enabled637d <= matchd636d;
	-- d638d
	sted638d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord638d,
			Enable=>Enabled638d,
			match=>matchd638d,
			run=>run);

	Enabled638d <= matchd637d;
	-- d639d
	sted639d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord639d,
			Enable=>Enabled639d,
			match=>matchd639d,
			run=>run);

	reports(24) <= matchd639d;
	Enabled639d <= matchd638d;
	-- d640d
	sted640d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord640d,
			Enable=>Enabled640d,
			match=>matchd640d,
			run=>run);

	-- d641d
	sted641d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord641d,
			Enable=>Enabled641d,
			match=>matchd641d,
			run=>run);

	Enabled641d <= matchd641d OR matchd640d;
	-- d642d
	sted642d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord642d,
			Enable=>Enabled642d,
			match=>matchd642d,
			run=>run);

	Enabled642d <= matchd641d;
	-- d643d
	sted643d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord643d,
			Enable=>Enabled643d,
			match=>matchd643d,
			run=>run);

	Enabled643d <= matchd642d;
	-- d644d
	sted644d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord644d,
			Enable=>Enabled644d,
			match=>matchd644d,
			run=>run);

	Enabled644d <= matchd643d;
	-- d645d
	sted645d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord645d,
			Enable=>Enabled645d,
			match=>matchd645d,
			run=>run);

	Enabled645d <= matchd644d;
	-- d646d
	sted646d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord646d,
			Enable=>Enabled646d,
			match=>matchd646d,
			run=>run);

	Enabled646d <= matchd645d;
	-- d647d
	sted647d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord647d,
			Enable=>Enabled647d,
			match=>matchd647d,
			run=>run);

	Enabled647d <= matchd646d OR matchd647d;
	-- d648d
	sted648d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord648d,
			Enable=>Enabled648d,
			match=>matchd648d,
			run=>run);

	Enabled648d <= matchd647d;
	-- d649d
	sted649d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord649d,
			Enable=>Enabled649d,
			match=>matchd649d,
			run=>run);

	Enabled649d <= matchd648d;
	-- d650d
	sted650d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord650d,
			Enable=>Enabled650d,
			match=>matchd650d,
			run=>run);

	Enabled650d <= matchd649d;
	-- d651d
	sted651d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord651d,
			Enable=>Enabled651d,
			match=>matchd651d,
			run=>run);

	reports(25) <= matchd651d;
	Enabled651d <= matchd650d;
	-- d652d
	sted652d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord652d,
			Enable=>Enabled652d,
			match=>matchd652d,
			run=>run);

	-- d653d
	sted653d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord653d,
			Enable=>Enabled653d,
			match=>matchd653d,
			run=>run);

	Enabled653d <= matchd653d OR matchd652d;
	-- d654d
	sted654d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord654d,
			Enable=>Enabled654d,
			match=>matchd654d,
			run=>run);

	Enabled654d <= matchd653d;
	-- d655d
	sted655d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord655d,
			Enable=>Enabled655d,
			match=>matchd655d,
			run=>run);

	Enabled655d <= matchd654d;
	-- d656d
	sted656d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord656d,
			Enable=>Enabled656d,
			match=>matchd656d,
			run=>run);

	Enabled656d <= matchd655d;
	-- d657d
	sted657d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord657d,
			Enable=>Enabled657d,
			match=>matchd657d,
			run=>run);

	Enabled657d <= matchd656d;
	-- d658d
	sted658d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord658d,
			Enable=>Enabled658d,
			match=>matchd658d,
			run=>run);

	Enabled658d <= matchd657d OR matchd658d;
	-- d659d
	sted659d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord659d,
			Enable=>Enabled659d,
			match=>matchd659d,
			run=>run);

	Enabled659d <= matchd658d;
	-- d660d
	sted660d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord660d,
			Enable=>Enabled660d,
			match=>matchd660d,
			run=>run);

	Enabled660d <= matchd659d;
	-- d661d
	sted661d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord661d,
			Enable=>Enabled661d,
			match=>matchd661d,
			run=>run);

	Enabled661d <= matchd660d;
	-- d662d
	sted662d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord662d,
			Enable=>Enabled662d,
			match=>matchd662d,
			run=>run);

	reports(26) <= matchd662d;
	Enabled662d <= matchd661d;
	-- d663d
	sted663d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord663d,
			Enable=>Enabled663d,
			match=>matchd663d,
			run=>run);

	-- d664d
	sted664d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord664d,
			Enable=>Enabled664d,
			match=>matchd664d,
			run=>run);

	Enabled664d <= matchd663d OR matchd664d;
	-- d665d
	sted665d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord665d,
			Enable=>Enabled665d,
			match=>matchd665d,
			run=>run);

	Enabled665d <= matchd664d;
	-- d666d
	sted666d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord666d,
			Enable=>Enabled666d,
			match=>matchd666d,
			run=>run);

	Enabled666d <= matchd665d;
	-- d667d
	sted667d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord667d,
			Enable=>Enabled667d,
			match=>matchd667d,
			run=>run);

	Enabled667d <= matchd666d;
	-- d668d
	sted668d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord668d,
			Enable=>Enabled668d,
			match=>matchd668d,
			run=>run);

	Enabled668d <= matchd667d;
	-- d669d
	sted669d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord669d,
			Enable=>Enabled669d,
			match=>matchd669d,
			run=>run);

	Enabled669d <= matchd668d OR matchd669d;
	-- d670d
	sted670d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord670d,
			Enable=>Enabled670d,
			match=>matchd670d,
			run=>run);

	Enabled670d <= matchd669d;
	-- d671d
	sted671d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord671d,
			Enable=>Enabled671d,
			match=>matchd671d,
			run=>run);

	Enabled671d <= matchd670d;
	-- d672d
	sted672d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord672d,
			Enable=>Enabled672d,
			match=>matchd672d,
			run=>run);

	Enabled672d <= matchd671d;
	-- d673d
	sted673d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord673d,
			Enable=>Enabled673d,
			match=>matchd673d,
			run=>run);

	Enabled673d <= matchd672d;
	-- d674d
	sted674d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord674d,
			Enable=>Enabled674d,
			match=>matchd674d,
			run=>run);

	reports(27) <= matchd674d;
	Enabled674d <= matchd673d;
	-- d675d
	sted675d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord675d,
			Enable=>Enabled675d,
			match=>matchd675d,
			run=>run);

	-- d676d
	sted676d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord676d,
			Enable=>Enabled676d,
			match=>matchd676d,
			run=>run);

	Enabled676d <= matchd676d OR matchd675d;
	-- d677d
	sted677d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord677d,
			Enable=>Enabled677d,
			match=>matchd677d,
			run=>run);

	Enabled677d <= matchd676d;
	-- d678d
	sted678d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord678d,
			Enable=>Enabled678d,
			match=>matchd678d,
			run=>run);

	Enabled678d <= matchd677d;
	-- d679d
	sted679d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord679d,
			Enable=>Enabled679d,
			match=>matchd679d,
			run=>run);

	Enabled679d <= matchd678d;
	-- d680d
	sted680d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord680d,
			Enable=>Enabled680d,
			match=>matchd680d,
			run=>run);

	Enabled680d <= matchd679d;
	-- d681d
	sted681d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord681d,
			Enable=>Enabled681d,
			match=>matchd681d,
			run=>run);

	Enabled681d <= matchd680d OR matchd681d;
	-- d682d
	sted682d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord682d,
			Enable=>Enabled682d,
			match=>matchd682d,
			run=>run);

	Enabled682d <= matchd681d;
	-- d683d
	sted683d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord683d,
			Enable=>Enabled683d,
			match=>matchd683d,
			run=>run);

	Enabled683d <= matchd682d;
	-- d684d
	sted684d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord684d,
			Enable=>Enabled684d,
			match=>matchd684d,
			run=>run);

	Enabled684d <= matchd683d;
	-- d685d
	sted685d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord685d,
			Enable=>Enabled685d,
			match=>matchd685d,
			run=>run);

	Enabled685d <= matchd684d;
	-- d686d
	sted686d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord686d,
			Enable=>Enabled686d,
			match=>matchd686d,
			run=>run);

	Enabled686d <= matchd686d OR matchd685d;
	-- d687d
	sted687d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord687d,
			Enable=>Enabled687d,
			match=>matchd687d,
			run=>run);

	Enabled687d <= matchd686d;
	-- d688d
	sted688d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord688d,
			Enable=>Enabled688d,
			match=>matchd688d,
			run=>run);

	Enabled688d <= matchd687d;
	-- d689d
	sted689d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord689d,
			Enable=>Enabled689d,
			match=>matchd689d,
			run=>run);

	Enabled689d <= matchd688d;
	-- d690d
	sted690d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord690d,
			Enable=>Enabled690d,
			match=>matchd690d,
			run=>run);

	reports(28) <= matchd690d;
	Enabled690d <= matchd689d;
	-- d691d
	sted691d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord691d,
			Enable=>Enabled691d,
			match=>matchd691d,
			run=>run);

	-- d692d
	sted692d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord692d,
			Enable=>Enabled692d,
			match=>matchd692d,
			run=>run);

	Enabled692d <= matchd691d OR matchd692d;
	-- d693d
	sted693d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord693d,
			Enable=>Enabled693d,
			match=>matchd693d,
			run=>run);

	Enabled693d <= matchd692d;
	-- d694d
	sted694d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord694d,
			Enable=>Enabled694d,
			match=>matchd694d,
			run=>run);

	Enabled694d <= matchd694d OR matchd693d;
	-- d695d
	sted695d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord695d,
			Enable=>Enabled695d,
			match=>matchd695d,
			run=>run);

	Enabled695d <= matchd694d;
	-- d696d
	sted696d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord696d,
			Enable=>Enabled696d,
			match=>matchd696d,
			run=>run);

	Enabled696d <= matchd695d OR matchd696d;
	-- d697d
	sted697d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord697d,
			Enable=>Enabled697d,
			match=>matchd697d,
			run=>run);

	Enabled697d <= matchd696d;
	-- d698d
	sted698d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord698d,
			Enable=>Enabled698d,
			match=>matchd698d,
			run=>run);

	Enabled698d <= matchd697d;
	-- d699d
	sted699d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord699d,
			Enable=>Enabled699d,
			match=>matchd699d,
			run=>run);

	Enabled699d <= matchd698d;
	-- d700d
	sted700d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord700d,
			Enable=>Enabled700d,
			match=>matchd700d,
			run=>run);

	Enabled700d <= matchd699d;
	-- d701d
	sted701d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord701d,
			Enable=>Enabled701d,
			match=>matchd701d,
			run=>run);

	Enabled701d <= matchd700d;
	-- d702d
	sted702d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord702d,
			Enable=>Enabled702d,
			match=>matchd702d,
			run=>run);

	Enabled702d <= matchd702d OR matchd701d;
	-- d703d
	sted703d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord703d,
			Enable=>Enabled703d,
			match=>matchd703d,
			run=>run);

	Enabled703d <= matchd702d;
	-- d704d
	sted704d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord704d,
			Enable=>Enabled704d,
			match=>matchd704d,
			run=>run);

	Enabled704d <= matchd703d;
	-- d705d
	sted705d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord705d,
			Enable=>Enabled705d,
			match=>matchd705d,
			run=>run);

	Enabled705d <= matchd704d;
	-- d706d
	sted706d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord706d,
			Enable=>Enabled706d,
			match=>matchd706d,
			run=>run);

	Enabled706d <= matchd705d;
	-- d707d
	sted707d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord707d,
			Enable=>Enabled707d,
			match=>matchd707d,
			run=>run);

	Enabled707d <= matchd706d;
	-- d708d
	sted708d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord708d,
			Enable=>Enabled708d,
			match=>matchd708d,
			run=>run);

	-- d709d
	sted709d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord709d,
			Enable=>Enabled709d,
			match=>matchd709d,
			run=>run);

	Enabled709d <= matchd709d OR matchd708d;
	-- d710d
	sted710d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord710d,
			Enable=>Enabled710d,
			match=>matchd710d,
			run=>run);

	Enabled710d <= matchd709d;
	-- d711d
	sted711d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord711d,
			Enable=>Enabled711d,
			match=>matchd711d,
			run=>run);

	Enabled711d <= matchd710d;
	-- d712d
	sted712d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord712d,
			Enable=>Enabled712d,
			match=>matchd712d,
			run=>run);

	Enabled712d <= matchd711d;
	-- d713d
	sted713d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord713d,
			Enable=>Enabled713d,
			match=>matchd713d,
			run=>run);

	Enabled713d <= matchd712d;
	-- d714d
	sted714d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord714d,
			Enable=>Enabled714d,
			match=>matchd714d,
			run=>run);

	Enabled714d <= matchd713d;
	-- d715d
	sted715d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord715d,
			Enable=>Enabled715d,
			match=>matchd715d,
			run=>run);

	Enabled715d <= matchd714d OR matchd715d;
	-- d716d
	sted716d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord716d,
			Enable=>Enabled716d,
			match=>matchd716d,
			run=>run);

	Enabled716d <= matchd715d;
	-- d717d
	sted717d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord717d,
			Enable=>Enabled717d,
			match=>matchd717d,
			run=>run);

	Enabled717d <= matchd716d OR matchd717d;
	-- d718d
	sted718d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord718d,
			Enable=>Enabled718d,
			match=>matchd718d,
			run=>run);

	Enabled718d <= matchd717d;
	-- d719d
	sted719d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord719d,
			Enable=>Enabled719d,
			match=>matchd719d,
			run=>run);

	Enabled719d <= matchd718d OR matchd719d;
	-- d720d
	sted720d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord720d,
			Enable=>Enabled720d,
			match=>matchd720d,
			run=>run);

	Enabled720d <= matchd719d;
	-- d721d
	sted721d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord721d,
			Enable=>Enabled721d,
			match=>matchd721d,
			run=>run);

	Enabled721d <= matchd720d;
	-- d722d
	sted722d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord722d,
			Enable=>Enabled722d,
			match=>matchd722d,
			run=>run);

	Enabled722d <= matchd721d;
	-- d723d
	sted723d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord723d,
			Enable=>Enabled723d,
			match=>matchd723d,
			run=>run);

	Enabled723d <= matchd722d;
	-- d724d
	sted724d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord724d,
			Enable=>Enabled724d,
			match=>matchd724d,
			run=>run);

	Enabled724d <= matchd723d;
	-- d726d
	sted726d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord726d,
			Enable=>Enabled726d,
			match=>matchd726d,
			run=>run);

	-- d727d
	sted727d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord727d,
			Enable=>Enabled727d,
			match=>matchd727d,
			run=>run);

	Enabled727d <= matchd727d OR matchd726d;
	-- d728d
	sted728d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord728d,
			Enable=>Enabled728d,
			match=>matchd728d,
			run=>run);

	Enabled728d <= matchd727d;
	-- d729d
	sted729d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord729d,
			Enable=>Enabled729d,
			match=>matchd729d,
			run=>run);

	Enabled729d <= matchd728d;
	-- d730d
	sted730d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord730d,
			Enable=>Enabled730d,
			match=>matchd730d,
			run=>run);

	Enabled730d <= matchd729d;
	-- d731d
	sted731d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord731d,
			Enable=>Enabled731d,
			match=>matchd731d,
			run=>run);

	Enabled731d <= matchd730d;
	-- d732d
	sted732d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord732d,
			Enable=>Enabled732d,
			match=>matchd732d,
			run=>run);

	Enabled732d <= matchd731d;
	-- d733d
	sted733d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord733d,
			Enable=>Enabled733d,
			match=>matchd733d,
			run=>run);

	Enabled733d <= matchd732d OR matchd733d;
	-- d734d
	sted734d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord734d,
			Enable=>Enabled734d,
			match=>matchd734d,
			run=>run);

	Enabled734d <= matchd733d;
	-- d735d
	sted735d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord735d,
			Enable=>Enabled735d,
			match=>matchd735d,
			run=>run);

	Enabled735d <= matchd734d;
	-- d736d
	sted736d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord736d,
			Enable=>Enabled736d,
			match=>matchd736d,
			run=>run);

	Enabled736d <= matchd735d;
	-- d737d
	sted737d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord737d,
			Enable=>Enabled737d,
			match=>matchd737d,
			run=>run);

	Enabled737d <= matchd736d;
	-- d738d
	sted738d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord738d,
			Enable=>Enabled738d,
			match=>matchd738d,
			run=>run);

	reports(29) <= matchd738d;
	Enabled738d <= matchd737d;
	-- d739d
	sted739d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord739d,
			Enable=>Enabled739d,
			match=>matchd739d,
			run=>run);

	-- d740d
	sted740d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord740d,
			Enable=>Enabled740d,
			match=>matchd740d,
			run=>run);

	Enabled740d <= matchd739d OR matchd740d;
	-- d741d
	sted741d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord741d,
			Enable=>Enabled741d,
			match=>matchd741d,
			run=>run);

	Enabled741d <= matchd740d;
	-- d742d
	sted742d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord742d,
			Enable=>Enabled742d,
			match=>matchd742d,
			run=>run);

	Enabled742d <= matchd741d;
	-- d743d
	sted743d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord743d,
			Enable=>Enabled743d,
			match=>matchd743d,
			run=>run);

	Enabled743d <= matchd742d;
	-- d744d
	sted744d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord744d,
			Enable=>Enabled744d,
			match=>matchd744d,
			run=>run);

	Enabled744d <= matchd743d;
	-- d745d
	sted745d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord745d,
			Enable=>Enabled745d,
			match=>matchd745d,
			run=>run);

	Enabled745d <= matchd745d OR matchd744d;
	-- d746d
	sted746d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord746d,
			Enable=>Enabled746d,
			match=>matchd746d,
			run=>run);

	Enabled746d <= matchd745d;
	-- d747d
	sted747d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord747d,
			Enable=>Enabled747d,
			match=>matchd747d,
			run=>run);

	Enabled747d <= matchd746d;
	-- d748d
	sted748d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord748d,
			Enable=>Enabled748d,
			match=>matchd748d,
			run=>run);

	Enabled748d <= matchd747d;
	-- d749d
	sted749d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord749d,
			Enable=>Enabled749d,
			match=>matchd749d,
			run=>run);

	Enabled749d <= matchd748d;
	-- d750d
	sted750d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord750d,
			Enable=>Enabled750d,
			match=>matchd750d,
			run=>run);

	reports(30) <= matchd750d;
	Enabled750d <= matchd749d;
	-- d751d
	sted751d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord751d,
			Enable=>Enabled751d,
			match=>matchd751d,
			run=>run);

	-- d752d
	sted752d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord752d,
			Enable=>Enabled752d,
			match=>matchd752d,
			run=>run);

	Enabled752d <= matchd751d;
	-- d753d
	sted753d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord753d,
			Enable=>Enabled753d,
			match=>matchd753d,
			run=>run);

	Enabled753d <= matchd752d;
	-- d754d
	sted754d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord754d,
			Enable=>Enabled754d,
			match=>matchd754d,
			run=>run);

	Enabled754d <= matchd753d;
	-- d755d
	sted755d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord755d,
			Enable=>Enabled755d,
			match=>matchd755d,
			run=>run);

	Enabled755d <= matchd754d;
	-- d756d
	sted756d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord756d,
			Enable=>Enabled756d,
			match=>matchd756d,
			run=>run);

	Enabled756d <= matchd755d;
	-- d757d
	sted757d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord757d,
			Enable=>Enabled757d,
			match=>matchd757d,
			run=>run);

	Enabled757d <= matchd756d;
	-- d758d
	sted758d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord758d,
			Enable=>Enabled758d,
			match=>matchd758d,
			run=>run);

	Enabled758d <= matchd757d;
	-- d759d
	sted759d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord759d,
			Enable=>Enabled759d,
			match=>matchd759d,
			run=>run);

	Enabled759d <= matchd758d;
	-- d760d
	sted760d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord760d,
			Enable=>Enabled760d,
			match=>matchd760d,
			run=>run);

	Enabled760d <= matchd759d;
	-- d761d
	sted761d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord761d,
			Enable=>Enabled761d,
			match=>matchd761d,
			run=>run);

	Enabled761d <= matchd761d OR matchd760d;
	-- d762d
	sted762d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord762d,
			Enable=>Enabled762d,
			match=>matchd762d,
			run=>run);

	Enabled762d <= matchd761d;
	-- d763d
	sted763d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord763d,
			Enable=>Enabled763d,
			match=>matchd763d,
			run=>run);

	Enabled763d <= matchd762d;
	-- d764d
	sted764d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord764d,
			Enable=>Enabled764d,
			match=>matchd764d,
			run=>run);

	Enabled764d <= matchd763d;
	-- d765d
	sted765d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord765d,
			Enable=>Enabled765d,
			match=>matchd765d,
			run=>run);

	reports(31) <= matchd765d;
	Enabled765d <= matchd764d;
	-- d766d
	sted766d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord766d,
			Enable=>Enabled766d,
			match=>matchd766d,
			run=>run);

	-- d767d
	sted767d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord767d,
			Enable=>Enabled767d,
			match=>matchd767d,
			run=>run);

	Enabled767d <= matchd767d OR matchd766d;
	-- d768d
	sted768d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord768d,
			Enable=>Enabled768d,
			match=>matchd768d,
			run=>run);

	Enabled768d <= matchd767d;
	-- d769d
	sted769d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord769d,
			Enable=>Enabled769d,
			match=>matchd769d,
			run=>run);

	Enabled769d <= matchd768d;
	-- d770d
	sted770d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord770d,
			Enable=>Enabled770d,
			match=>matchd770d,
			run=>run);

	Enabled770d <= matchd769d;
	-- d771d
	sted771d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord771d,
			Enable=>Enabled771d,
			match=>matchd771d,
			run=>run);

	Enabled771d <= matchd770d;
	-- d772d
	sted772d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord772d,
			Enable=>Enabled772d,
			match=>matchd772d,
			run=>run);

	Enabled772d <= matchd772d OR matchd771d;
	-- d773d
	sted773d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord773d,
			Enable=>Enabled773d,
			match=>matchd773d,
			run=>run);

	Enabled773d <= matchd772d;
	-- d774d
	sted774d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord774d,
			Enable=>Enabled774d,
			match=>matchd774d,
			run=>run);

	Enabled774d <= matchd773d;
	-- d775d
	sted775d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord775d,
			Enable=>Enabled775d,
			match=>matchd775d,
			run=>run);

	Enabled775d <= matchd774d;
	-- d776d
	sted776d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord776d,
			Enable=>Enabled776d,
			match=>matchd776d,
			run=>run);

	reports(32) <= matchd776d;
	Enabled776d <= matchd775d;
	-- d777d
	sted777d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord777d,
			Enable=>Enabled777d,
			match=>matchd777d,
			run=>run);

	-- d778d
	sted778d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord778d,
			Enable=>Enabled778d,
			match=>matchd778d,
			run=>run);

	Enabled778d <= matchd777d OR matchd778d;
	-- d779d
	sted779d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord779d,
			Enable=>Enabled779d,
			match=>matchd779d,
			run=>run);

	Enabled779d <= matchd778d;
	-- d780d
	sted780d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord780d,
			Enable=>Enabled780d,
			match=>matchd780d,
			run=>run);

	Enabled780d <= matchd779d;
	-- d781d
	sted781d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord781d,
			Enable=>Enabled781d,
			match=>matchd781d,
			run=>run);

	Enabled781d <= matchd780d;
	-- d782d
	sted782d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord782d,
			Enable=>Enabled782d,
			match=>matchd782d,
			run=>run);

	Enabled782d <= matchd781d;
	-- d783d
	sted783d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord783d,
			Enable=>Enabled783d,
			match=>matchd783d,
			run=>run);

	Enabled783d <= matchd783d OR matchd782d;
	-- d784d
	sted784d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord784d,
			Enable=>Enabled784d,
			match=>matchd784d,
			run=>run);

	Enabled784d <= matchd783d;
	-- d785d
	sted785d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord785d,
			Enable=>Enabled785d,
			match=>matchd785d,
			run=>run);

	Enabled785d <= matchd784d;
	-- d786d
	sted786d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord786d,
			Enable=>Enabled786d,
			match=>matchd786d,
			run=>run);

	Enabled786d <= matchd785d;
	-- d787d
	sted787d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord787d,
			Enable=>Enabled787d,
			match=>matchd787d,
			run=>run);

	reports(33) <= matchd787d;
	Enabled787d <= matchd786d;
	-- d788d
	sted788d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord788d,
			Enable=>Enabled788d,
			match=>matchd788d,
			run=>run);

	-- d789d
	sted789d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord789d,
			Enable=>Enabled789d,
			match=>matchd789d,
			run=>run);

	Enabled789d <= matchd789d OR matchd788d;
	-- d790d
	sted790d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord790d,
			Enable=>Enabled790d,
			match=>matchd790d,
			run=>run);

	Enabled790d <= matchd789d;
	-- d791d
	sted791d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord791d,
			Enable=>Enabled791d,
			match=>matchd791d,
			run=>run);

	Enabled791d <= matchd790d;
	-- d792d
	sted792d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord792d,
			Enable=>Enabled792d,
			match=>matchd792d,
			run=>run);

	Enabled792d <= matchd791d;
	-- d793d
	sted793d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord793d,
			Enable=>Enabled793d,
			match=>matchd793d,
			run=>run);

	Enabled793d <= matchd792d;
	-- d794d
	sted794d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord794d,
			Enable=>Enabled794d,
			match=>matchd794d,
			run=>run);

	Enabled794d <= matchd793d OR matchd794d;
	-- d795d
	sted795d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord795d,
			Enable=>Enabled795d,
			match=>matchd795d,
			run=>run);

	Enabled795d <= matchd794d;
	-- d796d
	sted796d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord796d,
			Enable=>Enabled796d,
			match=>matchd796d,
			run=>run);

	Enabled796d <= matchd795d;
	-- d797d
	sted797d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord797d,
			Enable=>Enabled797d,
			match=>matchd797d,
			run=>run);

	Enabled797d <= matchd796d;
	-- d798d
	sted798d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord798d,
			Enable=>Enabled798d,
			match=>matchd798d,
			run=>run);

	Enabled798d <= matchd797d;
	-- d799d
	sted799d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord799d,
			Enable=>Enabled799d,
			match=>matchd799d,
			run=>run);

	Enabled799d <= matchd798d OR matchd799d;
	-- d800d
	sted800d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord800d,
			Enable=>Enabled800d,
			match=>matchd800d,
			run=>run);

	Enabled800d <= matchd799d;
	-- d801d
	sted801d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord801d,
			Enable=>Enabled801d,
			match=>matchd801d,
			run=>run);

	Enabled801d <= matchd801d OR matchd800d;
	-- d802d
	sted802d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord802d,
			Enable=>Enabled802d,
			match=>matchd802d,
			run=>run);

	Enabled802d <= matchd801d;
	-- d803d
	sted803d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord803d,
			Enable=>Enabled803d,
			match=>matchd803d,
			run=>run);

	-- d804d
	sted804d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord804d,
			Enable=>Enabled804d,
			match=>matchd804d,
			run=>run);

	Enabled804d <= matchd803d OR matchd804d;
	-- d805d
	sted805d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord805d,
			Enable=>Enabled805d,
			match=>matchd805d,
			run=>run);

	Enabled805d <= matchd804d;
	-- d806d
	sted806d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord806d,
			Enable=>Enabled806d,
			match=>matchd806d,
			run=>run);

	Enabled806d <= matchd805d;
	-- d807d
	sted807d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord807d,
			Enable=>Enabled807d,
			match=>matchd807d,
			run=>run);

	Enabled807d <= matchd806d;
	-- d808d
	sted808d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord808d,
			Enable=>Enabled808d,
			match=>matchd808d,
			run=>run);

	Enabled808d <= matchd807d;
	-- d809d
	sted809d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord809d,
			Enable=>Enabled809d,
			match=>matchd809d,
			run=>run);

	Enabled809d <= matchd808d OR matchd809d;
	-- d810d
	sted810d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord810d,
			Enable=>Enabled810d,
			match=>matchd810d,
			run=>run);

	Enabled810d <= matchd809d;
	-- d811d
	sted811d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord811d,
			Enable=>Enabled811d,
			match=>matchd811d,
			run=>run);

	Enabled811d <= matchd811d OR matchd810d;
	-- d812d
	sted812d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord812d,
			Enable=>Enabled812d,
			match=>matchd812d,
			run=>run);

	Enabled812d <= matchd811d;
	-- d813d
	sted813d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord813d,
			Enable=>Enabled813d,
			match=>matchd813d,
			run=>run);

	Enabled813d <= matchd813d OR matchd812d;
	-- d814d
	sted814d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord814d,
			Enable=>Enabled814d,
			match=>matchd814d,
			run=>run);

	Enabled814d <= matchd813d;
	-- d815d
	sted815d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord815d,
			Enable=>Enabled815d,
			match=>matchd815d,
			run=>run);

	Enabled815d <= matchd814d;
	-- d816d
	sted816d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord816d,
			Enable=>Enabled816d,
			match=>matchd816d,
			run=>run);

	Enabled816d <= matchd815d;
	-- d817d
	sted817d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord817d,
			Enable=>Enabled817d,
			match=>matchd817d,
			run=>run);

	Enabled817d <= matchd816d;
	-- d819d
	sted819d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord819d,
			Enable=>Enabled819d,
			match=>matchd819d,
			run=>run);

	-- d820d
	sted820d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord820d,
			Enable=>Enabled820d,
			match=>matchd820d,
			run=>run);

	Enabled820d <= matchd819d OR matchd820d;
	-- d821d
	sted821d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord821d,
			Enable=>Enabled821d,
			match=>matchd821d,
			run=>run);

	Enabled821d <= matchd820d;
	-- d822d
	sted822d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord822d,
			Enable=>Enabled822d,
			match=>matchd822d,
			run=>run);

	Enabled822d <= matchd821d;
	-- d823d
	sted823d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord823d,
			Enable=>Enabled823d,
			match=>matchd823d,
			run=>run);

	Enabled823d <= matchd822d;
	-- d824d
	sted824d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord824d,
			Enable=>Enabled824d,
			match=>matchd824d,
			run=>run);

	Enabled824d <= matchd823d;
	-- d825d
	sted825d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord825d,
			Enable=>Enabled825d,
			match=>matchd825d,
			run=>run);

	Enabled825d <= matchd824d;
	-- d826d
	sted826d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord826d,
			Enable=>Enabled826d,
			match=>matchd826d,
			run=>run);

	Enabled826d <= matchd825d OR matchd826d;
	-- d827d
	sted827d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord827d,
			Enable=>Enabled827d,
			match=>matchd827d,
			run=>run);

	Enabled827d <= matchd826d;
	-- d828d
	sted828d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord828d,
			Enable=>Enabled828d,
			match=>matchd828d,
			run=>run);

	Enabled828d <= matchd827d;
	-- d829d
	sted829d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord829d,
			Enable=>Enabled829d,
			match=>matchd829d,
			run=>run);

	Enabled829d <= matchd828d;
	-- d830d
	sted830d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord830d,
			Enable=>Enabled830d,
			match=>matchd830d,
			run=>run);

	reports(34) <= matchd830d;
	Enabled830d <= matchd829d;
	-- d831d
	sted831d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord831d,
			Enable=>Enabled831d,
			match=>matchd831d,
			run=>run);

	-- d832d
	sted832d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord832d,
			Enable=>Enabled832d,
			match=>matchd832d,
			run=>run);

	Enabled832d <= matchd831d OR matchd832d;
	-- d833d
	sted833d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord833d,
			Enable=>Enabled833d,
			match=>matchd833d,
			run=>run);

	Enabled833d <= matchd832d;
	-- d834d
	sted834d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord834d,
			Enable=>Enabled834d,
			match=>matchd834d,
			run=>run);

	Enabled834d <= matchd833d;
	-- d835d
	sted835d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord835d,
			Enable=>Enabled835d,
			match=>matchd835d,
			run=>run);

	Enabled835d <= matchd834d;
	-- d836d
	sted836d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord836d,
			Enable=>Enabled836d,
			match=>matchd836d,
			run=>run);

	Enabled836d <= matchd835d;
	-- d837d
	sted837d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord837d,
			Enable=>Enabled837d,
			match=>matchd837d,
			run=>run);

	Enabled837d <= matchd836d;
	-- d838d
	sted838d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord838d,
			Enable=>Enabled838d,
			match=>matchd838d,
			run=>run);

	Enabled838d <= matchd838d OR matchd837d;
	-- d839d
	sted839d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord839d,
			Enable=>Enabled839d,
			match=>matchd839d,
			run=>run);

	Enabled839d <= matchd838d;
	-- d840d
	sted840d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord840d,
			Enable=>Enabled840d,
			match=>matchd840d,
			run=>run);

	Enabled840d <= matchd839d;
	-- d841d
	sted841d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord841d,
			Enable=>Enabled841d,
			match=>matchd841d,
			run=>run);

	Enabled841d <= matchd840d;
	-- d842d
	sted842d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord842d,
			Enable=>Enabled842d,
			match=>matchd842d,
			run=>run);

	reports(35) <= matchd842d;
	Enabled842d <= matchd841d;
	-- d843d
	sted843d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord843d,
			Enable=>Enabled843d,
			match=>matchd843d,
			run=>run);

	-- d844d
	sted844d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord844d,
			Enable=>Enabled844d,
			match=>matchd844d,
			run=>run);

	Enabled844d <= matchd843d OR matchd844d;
	-- d845d
	sted845d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord845d,
			Enable=>Enabled845d,
			match=>matchd845d,
			run=>run);

	Enabled845d <= matchd844d;
	-- d846d
	sted846d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord846d,
			Enable=>Enabled846d,
			match=>matchd846d,
			run=>run);

	Enabled846d <= matchd845d;
	-- d847d
	sted847d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord847d,
			Enable=>Enabled847d,
			match=>matchd847d,
			run=>run);

	Enabled847d <= matchd846d;
	-- d848d
	sted848d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord848d,
			Enable=>Enabled848d,
			match=>matchd848d,
			run=>run);

	Enabled848d <= matchd847d;
	-- d849d
	sted849d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord849d,
			Enable=>Enabled849d,
			match=>matchd849d,
			run=>run);

	Enabled849d <= matchd848d;
	-- d850d
	sted850d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord850d,
			Enable=>Enabled850d,
			match=>matchd850d,
			run=>run);

	Enabled850d <= matchd849d OR matchd850d;
	-- d851d
	sted851d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord851d,
			Enable=>Enabled851d,
			match=>matchd851d,
			run=>run);

	Enabled851d <= matchd850d;
	-- d852d
	sted852d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord852d,
			Enable=>Enabled852d,
			match=>matchd852d,
			run=>run);

	Enabled852d <= matchd852d OR matchd851d;
	-- d853d
	sted853d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord853d,
			Enable=>Enabled853d,
			match=>matchd853d,
			run=>run);

	Enabled853d <= matchd852d;
	-- d854d
	sted854d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord854d,
			Enable=>Enabled854d,
			match=>matchd854d,
			run=>run);

	Enabled854d <= matchd853d OR matchd854d;
	-- d855d
	sted855d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord855d,
			Enable=>Enabled855d,
			match=>matchd855d,
			run=>run);

	Enabled855d <= matchd854d;
	-- d856d
	sted856d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord856d,
			Enable=>Enabled856d,
			match=>matchd856d,
			run=>run);

	Enabled856d <= matchd856d OR matchd855d;
	-- d857d
	sted857d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord857d,
			Enable=>Enabled857d,
			match=>matchd857d,
			run=>run);

	Enabled857d <= matchd856d;
	-- d858d
	sted858d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord858d,
			Enable=>Enabled858d,
			match=>matchd858d,
			run=>run);

	Enabled858d <= matchd857d OR matchd858d;
	-- d859d
	sted859d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord859d,
			Enable=>Enabled859d,
			match=>matchd859d,
			run=>run);

	Enabled859d <= matchd858d;
	-- d860d
	sted860d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord860d,
			Enable=>Enabled860d,
			match=>matchd860d,
			run=>run);

	Enabled860d <= matchd859d;
	-- d861d
	sted861d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord861d,
			Enable=>Enabled861d,
			match=>matchd861d,
			run=>run);

	Enabled861d <= matchd860d;
	-- d862d
	sted862d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord862d,
			Enable=>Enabled862d,
			match=>matchd862d,
			run=>run);

	Enabled862d <= matchd861d;
	-- d863d
	sted863d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord863d,
			Enable=>Enabled863d,
			match=>matchd863d,
			run=>run);

	Enabled863d <= matchd862d;
	-- d864d
	sted864d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord864d,
			Enable=>Enabled864d,
			match=>matchd864d,
			run=>run);

	-- d865d
	sted865d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord865d,
			Enable=>Enabled865d,
			match=>matchd865d,
			run=>run);

	Enabled865d <= matchd864d OR matchd865d;
	-- d866d
	sted866d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord866d,
			Enable=>Enabled866d,
			match=>matchd866d,
			run=>run);

	Enabled866d <= matchd865d;
	-- d867d
	sted867d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord867d,
			Enable=>Enabled867d,
			match=>matchd867d,
			run=>run);

	Enabled867d <= matchd867d OR matchd866d;
	-- d868d
	sted868d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord868d,
			Enable=>Enabled868d,
			match=>matchd868d,
			run=>run);

	Enabled868d <= matchd867d;
	-- d869d
	sted869d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord869d,
			Enable=>Enabled869d,
			match=>matchd869d,
			run=>run);

	Enabled869d <= matchd868d OR matchd869d;
	-- d870d
	sted870d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord870d,
			Enable=>Enabled870d,
			match=>matchd870d,
			run=>run);

	Enabled870d <= matchd869d;
	-- d871d
	sted871d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord871d,
			Enable=>Enabled871d,
			match=>matchd871d,
			run=>run);

	Enabled871d <= matchd870d;
	-- d872d
	sted872d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord872d,
			Enable=>Enabled872d,
			match=>matchd872d,
			run=>run);

	Enabled872d <= matchd871d;
	-- d873d
	sted873d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord873d,
			Enable=>Enabled873d,
			match=>matchd873d,
			run=>run);

	Enabled873d <= matchd872d;
	-- d874d
	sted874d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord874d,
			Enable=>Enabled874d,
			match=>matchd874d,
			run=>run);

	Enabled874d <= matchd873d;
	-- d875d
	sted875d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord875d,
			Enable=>Enabled875d,
			match=>matchd875d,
			run=>run);

	Enabled875d <= matchd875d OR matchd874d;
	-- d876d
	sted876d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord876d,
			Enable=>Enabled876d,
			match=>matchd876d,
			run=>run);

	Enabled876d <= matchd875d;
	-- d877d
	sted877d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord877d,
			Enable=>Enabled877d,
			match=>matchd877d,
			run=>run);

	Enabled877d <= matchd877d OR matchd876d;
	-- d878d
	sted878d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord878d,
			Enable=>Enabled878d,
			match=>matchd878d,
			run=>run);

	Enabled878d <= matchd877d;
	-- d879d
	sted879d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord879d,
			Enable=>Enabled879d,
			match=>matchd879d,
			run=>run);

	Enabled879d <= matchd879d OR matchd878d;
	-- d880d
	sted880d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord880d,
			Enable=>Enabled880d,
			match=>matchd880d,
			run=>run);

	Enabled880d <= matchd879d;
	-- d881d
	sted881d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord881d,
			Enable=>Enabled881d,
			match=>matchd881d,
			run=>run);

	Enabled881d <= matchd880d;
	-- d882d
	sted882d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord882d,
			Enable=>Enabled882d,
			match=>matchd882d,
			run=>run);

	Enabled882d <= matchd881d;
	-- d883d
	sted883d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord883d,
			Enable=>Enabled883d,
			match=>matchd883d,
			run=>run);

	Enabled883d <= matchd882d;
	-- d884d
	sted884d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord884d,
			Enable=>Enabled884d,
			match=>matchd884d,
			run=>run);

	Enabled884d <= matchd883d;
	-- d885d
	sted885d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord885d,
			Enable=>Enabled885d,
			match=>matchd885d,
			run=>run);

	-- d886d
	sted886d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord886d,
			Enable=>Enabled886d,
			match=>matchd886d,
			run=>run);

	Enabled886d <= matchd885d OR matchd886d;
	-- d887d
	sted887d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord887d,
			Enable=>Enabled887d,
			match=>matchd887d,
			run=>run);

	Enabled887d <= matchd886d;
	-- d888d
	sted888d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord888d,
			Enable=>Enabled888d,
			match=>matchd888d,
			run=>run);

	Enabled888d <= matchd887d OR matchd888d;
	-- d889d
	sted889d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord889d,
			Enable=>Enabled889d,
			match=>matchd889d,
			run=>run);

	Enabled889d <= matchd888d;
	-- d890d
	sted890d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord890d,
			Enable=>Enabled890d,
			match=>matchd890d,
			run=>run);

	Enabled890d <= matchd890d OR matchd889d;
	-- d891d
	sted891d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord891d,
			Enable=>Enabled891d,
			match=>matchd891d,
			run=>run);

	Enabled891d <= matchd890d;
	-- d892d
	sted892d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord892d,
			Enable=>Enabled892d,
			match=>matchd892d,
			run=>run);

	Enabled892d <= matchd892d OR matchd891d;
	-- d893d
	sted893d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord893d,
			Enable=>Enabled893d,
			match=>matchd893d,
			run=>run);

	Enabled893d <= matchd892d;
	-- d894d
	sted894d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord894d,
			Enable=>Enabled894d,
			match=>matchd894d,
			run=>run);

	Enabled894d <= matchd894d OR matchd893d;
	-- d895d
	sted895d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord895d,
			Enable=>Enabled895d,
			match=>matchd895d,
			run=>run);

	Enabled895d <= matchd894d;
	-- d896d
	sted896d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord896d,
			Enable=>Enabled896d,
			match=>matchd896d,
			run=>run);

	Enabled896d <= matchd895d;
	-- d897d
	sted897d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord897d,
			Enable=>Enabled897d,
			match=>matchd897d,
			run=>run);

	Enabled897d <= matchd896d;
	-- d898d
	sted898d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord898d,
			Enable=>Enabled898d,
			match=>matchd898d,
			run=>run);

	Enabled898d <= matchd897d;
	-- d899d
	sted899d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord899d,
			Enable=>Enabled899d,
			match=>matchd899d,
			run=>run);

	Enabled899d <= matchd898d;
	-- d900d
	sted900d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord900d,
			Enable=>Enabled900d,
			match=>matchd900d,
			run=>run);

	Enabled900d <= matchd900d OR matchd899d;
	-- d901d
	sted901d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord901d,
			Enable=>Enabled901d,
			match=>matchd901d,
			run=>run);

	Enabled901d <= matchd900d;
	-- d902d
	sted902d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord902d,
			Enable=>Enabled902d,
			match=>matchd902d,
			run=>run);

	Enabled902d <= matchd901d;
	-- d903d
	sted903d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord903d,
			Enable=>Enabled903d,
			match=>matchd903d,
			run=>run);

	Enabled903d <= matchd902d;
	-- d904d
	sted904d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord904d,
			Enable=>Enabled904d,
			match=>matchd904d,
			run=>run);

	Enabled904d <= matchd903d;
	-- d905d
	sted905d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord905d,
			Enable=>Enabled905d,
			match=>matchd905d,
			run=>run);

	Enabled905d <= matchd904d;
	-- d907d
	sted907d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord907d,
			Enable=>Enabled907d,
			match=>matchd907d,
			run=>run);

	-- d908d
	sted908d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord908d,
			Enable=>Enabled908d,
			match=>matchd908d,
			run=>run);

	Enabled908d <= matchd907d OR matchd908d;
	-- d909d
	sted909d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord909d,
			Enable=>Enabled909d,
			match=>matchd909d,
			run=>run);

	Enabled909d <= matchd908d;
	-- d910d
	sted910d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord910d,
			Enable=>Enabled910d,
			match=>matchd910d,
			run=>run);

	Enabled910d <= matchd909d;
	-- d911d
	sted911d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord911d,
			Enable=>Enabled911d,
			match=>matchd911d,
			run=>run);

	Enabled911d <= matchd910d;
	-- d912d
	sted912d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord912d,
			Enable=>Enabled912d,
			match=>matchd912d,
			run=>run);

	Enabled912d <= matchd911d;
	-- d913d
	sted913d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord913d,
			Enable=>Enabled913d,
			match=>matchd913d,
			run=>run);

	Enabled913d <= matchd912d;
	-- d914d
	sted914d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord914d,
			Enable=>Enabled914d,
			match=>matchd914d,
			run=>run);

	Enabled914d <= matchd913d OR matchd914d;
	-- d915d
	sted915d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord915d,
			Enable=>Enabled915d,
			match=>matchd915d,
			run=>run);

	Enabled915d <= matchd914d;
	-- d916d
	sted916d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord916d,
			Enable=>Enabled916d,
			match=>matchd916d,
			run=>run);

	Enabled916d <= matchd915d;
	-- d917d
	sted917d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord917d,
			Enable=>Enabled917d,
			match=>matchd917d,
			run=>run);

	Enabled917d <= matchd916d;
	-- d918d
	sted918d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord918d,
			Enable=>Enabled918d,
			match=>matchd918d,
			run=>run);

	reports(36) <= matchd918d;
	Enabled918d <= matchd917d;
	-- d919d
	sted919d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord919d,
			Enable=>Enabled919d,
			match=>matchd919d,
			run=>run);

	-- d920d
	sted920d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord920d,
			Enable=>Enabled920d,
			match=>matchd920d,
			run=>run);

	Enabled920d <= matchd920d OR matchd919d;
	-- d921d
	sted921d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord921d,
			Enable=>Enabled921d,
			match=>matchd921d,
			run=>run);

	Enabled921d <= matchd920d;
	-- d922d
	sted922d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord922d,
			Enable=>Enabled922d,
			match=>matchd922d,
			run=>run);

	Enabled922d <= matchd921d;
	-- d923d
	sted923d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord923d,
			Enable=>Enabled923d,
			match=>matchd923d,
			run=>run);

	Enabled923d <= matchd922d;
	-- d924d
	sted924d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord924d,
			Enable=>Enabled924d,
			match=>matchd924d,
			run=>run);

	Enabled924d <= matchd923d;
	-- d925d
	sted925d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord925d,
			Enable=>Enabled925d,
			match=>matchd925d,
			run=>run);

	Enabled925d <= matchd925d OR matchd924d;
	-- d926d
	sted926d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord926d,
			Enable=>Enabled926d,
			match=>matchd926d,
			run=>run);

	Enabled926d <= matchd925d;
	-- d927d
	sted927d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord927d,
			Enable=>Enabled927d,
			match=>matchd927d,
			run=>run);

	Enabled927d <= matchd926d;
	-- d928d
	sted928d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord928d,
			Enable=>Enabled928d,
			match=>matchd928d,
			run=>run);

	Enabled928d <= matchd927d;
	-- d929d
	sted929d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord929d,
			Enable=>Enabled929d,
			match=>matchd929d,
			run=>run);

	Enabled929d <= matchd928d;
	-- d930d
	sted930d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord930d,
			Enable=>Enabled930d,
			match=>matchd930d,
			run=>run);

	reports(37) <= matchd930d;
	Enabled930d <= matchd929d;
	-- d931d
	sted931d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord931d,
			Enable=>Enabled931d,
			match=>matchd931d,
			run=>run);

	-- d932d
	sted932d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord932d,
			Enable=>Enabled932d,
			match=>matchd932d,
			run=>run);

	Enabled932d <= matchd931d OR matchd932d;
	-- d933d
	sted933d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord933d,
			Enable=>Enabled933d,
			match=>matchd933d,
			run=>run);

	Enabled933d <= matchd932d;
	-- d934d
	sted934d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord934d,
			Enable=>Enabled934d,
			match=>matchd934d,
			run=>run);

	Enabled934d <= matchd933d;
	-- d935d
	sted935d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord935d,
			Enable=>Enabled935d,
			match=>matchd935d,
			run=>run);

	Enabled935d <= matchd934d;
	-- d936d
	sted936d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord936d,
			Enable=>Enabled936d,
			match=>matchd936d,
			run=>run);

	Enabled936d <= matchd935d;
	-- d937d
	sted937d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord937d,
			Enable=>Enabled937d,
			match=>matchd937d,
			run=>run);

	Enabled937d <= matchd936d;
	-- d938d
	sted938d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord938d,
			Enable=>Enabled938d,
			match=>matchd938d,
			run=>run);

	Enabled938d <= matchd938d OR matchd937d;
	-- d939d
	sted939d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord939d,
			Enable=>Enabled939d,
			match=>matchd939d,
			run=>run);

	Enabled939d <= matchd938d;
	-- d940d
	sted940d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord940d,
			Enable=>Enabled940d,
			match=>matchd940d,
			run=>run);

	Enabled940d <= matchd939d;
	-- d941d
	sted941d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord941d,
			Enable=>Enabled941d,
			match=>matchd941d,
			run=>run);

	Enabled941d <= matchd940d;
	-- d942d
	sted942d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord942d,
			Enable=>Enabled942d,
			match=>matchd942d,
			run=>run);

	reports(38) <= matchd942d;
	Enabled942d <= matchd941d;
	-- d943d
	sted943d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord943d,
			Enable=>Enabled943d,
			match=>matchd943d,
			run=>run);

	-- d944d
	sted944d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord944d,
			Enable=>Enabled944d,
			match=>matchd944d,
			run=>run);

	Enabled944d <= matchd943d;
	-- d945d
	sted945d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord945d,
			Enable=>Enabled945d,
			match=>matchd945d,
			run=>run);

	Enabled945d <= matchd944d;
	-- d946d
	sted946d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord946d,
			Enable=>Enabled946d,
			match=>matchd946d,
			run=>run);

	Enabled946d <= matchd945d;
	-- d947d
	sted947d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord947d,
			Enable=>Enabled947d,
			match=>matchd947d,
			run=>run);

	Enabled947d <= matchd946d;
	-- d948d
	sted948d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord948d,
			Enable=>Enabled948d,
			match=>matchd948d,
			run=>run);

	Enabled948d <= matchd947d;
	-- d949d
	sted949d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord949d,
			Enable=>Enabled949d,
			match=>matchd949d,
			run=>run);

	Enabled949d <= matchd948d;
	-- d950d
	sted950d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord950d,
			Enable=>Enabled950d,
			match=>matchd950d,
			run=>run);

	Enabled950d <= matchd949d;
	-- d951d
	sted951d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord951d,
			Enable=>Enabled951d,
			match=>matchd951d,
			run=>run);

	Enabled951d <= matchd950d;
	-- d952d
	sted952d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord952d,
			Enable=>Enabled952d,
			match=>matchd952d,
			run=>run);

	Enabled952d <= matchd951d;
	-- d953d
	sted953d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord953d,
			Enable=>Enabled953d,
			match=>matchd953d,
			run=>run);

	Enabled953d <= matchd952d OR matchd953d;
	-- d954d
	sted954d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord954d,
			Enable=>Enabled954d,
			match=>matchd954d,
			run=>run);

	Enabled954d <= matchd953d;
	-- d955d
	sted955d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord955d,
			Enable=>Enabled955d,
			match=>matchd955d,
			run=>run);

	Enabled955d <= matchd954d;
	-- d956d
	sted956d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord956d,
			Enable=>Enabled956d,
			match=>matchd956d,
			run=>run);

	reports(39) <= matchd956d;
	Enabled956d <= matchd955d;
	-- d957d
	sted957d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord957d,
			Enable=>Enabled957d,
			match=>matchd957d,
			run=>run);

	-- d958d
	sted958d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord958d,
			Enable=>Enabled958d,
			match=>matchd958d,
			run=>run);

	Enabled958d <= matchd958d OR matchd957d;
	-- d959d
	sted959d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord959d,
			Enable=>Enabled959d,
			match=>matchd959d,
			run=>run);

	Enabled959d <= matchd958d;
	-- d960d
	sted960d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord960d,
			Enable=>Enabled960d,
			match=>matchd960d,
			run=>run);

	Enabled960d <= matchd959d;
	-- d961d
	sted961d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord961d,
			Enable=>Enabled961d,
			match=>matchd961d,
			run=>run);

	Enabled961d <= matchd960d;
	-- d962d
	sted962d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord962d,
			Enable=>Enabled962d,
			match=>matchd962d,
			run=>run);

	Enabled962d <= matchd961d;
	-- d963d
	sted963d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord963d,
			Enable=>Enabled963d,
			match=>matchd963d,
			run=>run);

	Enabled963d <= matchd963d OR matchd962d;
	-- d964d
	sted964d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord964d,
			Enable=>Enabled964d,
			match=>matchd964d,
			run=>run);

	Enabled964d <= matchd963d;
	-- d965d
	sted965d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord965d,
			Enable=>Enabled965d,
			match=>matchd965d,
			run=>run);

	Enabled965d <= matchd964d;
	-- d966d
	sted966d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord966d,
			Enable=>Enabled966d,
			match=>matchd966d,
			run=>run);

	Enabled966d <= matchd965d;
	-- d967d
	sted967d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord967d,
			Enable=>Enabled967d,
			match=>matchd967d,
			run=>run);

	Enabled967d <= matchd967d OR matchd966d;
	-- d968d
	sted968d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord968d,
			Enable=>Enabled968d,
			match=>matchd968d,
			run=>run);

	Enabled968d <= matchd967d;
	-- d969d
	sted969d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord969d,
			Enable=>Enabled969d,
			match=>matchd969d,
			run=>run);

	Enabled969d <= matchd969d OR matchd968d;
	-- d970d
	sted970d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord970d,
			Enable=>Enabled970d,
			match=>matchd970d,
			run=>run);

	Enabled970d <= matchd969d;
	-- d971d
	sted971d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord971d,
			Enable=>Enabled971d,
			match=>matchd971d,
			run=>run);

	-- d972d
	sted972d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord972d,
			Enable=>Enabled972d,
			match=>matchd972d,
			run=>run);

	Enabled972d <= matchd971d OR matchd972d;
	-- d973d
	sted973d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord973d,
			Enable=>Enabled973d,
			match=>matchd973d,
			run=>run);

	Enabled973d <= matchd972d;
	-- d974d
	sted974d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord974d,
			Enable=>Enabled974d,
			match=>matchd974d,
			run=>run);

	Enabled974d <= matchd973d;
	-- d975d
	sted975d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord975d,
			Enable=>Enabled975d,
			match=>matchd975d,
			run=>run);

	Enabled975d <= matchd974d;
	-- d976d
	sted976d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord976d,
			Enable=>Enabled976d,
			match=>matchd976d,
			run=>run);

	Enabled976d <= matchd975d;
	-- d977d
	sted977d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord977d,
			Enable=>Enabled977d,
			match=>matchd977d,
			run=>run);

	Enabled977d <= matchd976d OR matchd977d;
	-- d978d
	sted978d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord978d,
			Enable=>Enabled978d,
			match=>matchd978d,
			run=>run);

	Enabled978d <= matchd977d;
	-- d979d
	sted979d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord979d,
			Enable=>Enabled979d,
			match=>matchd979d,
			run=>run);

	Enabled979d <= matchd978d OR matchd979d;
	-- d980d
	sted980d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord980d,
			Enable=>Enabled980d,
			match=>matchd980d,
			run=>run);

	Enabled980d <= matchd979d;
	-- d981d
	sted981d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord981d,
			Enable=>Enabled981d,
			match=>matchd981d,
			run=>run);

	Enabled981d <= matchd981d OR matchd980d;
	-- d982d
	sted982d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord982d,
			Enable=>Enabled982d,
			match=>matchd982d,
			run=>run);

	Enabled982d <= matchd981d;
	-- d983d
	sted983d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord983d,
			Enable=>Enabled983d,
			match=>matchd983d,
			run=>run);

	Enabled983d <= matchd982d;
	-- d984d
	sted984d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord984d,
			Enable=>Enabled984d,
			match=>matchd984d,
			run=>run);

	Enabled984d <= matchd983d;
	-- d986d
	sted986d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord986d,
			Enable=>Enabled986d,
			match=>matchd986d,
			run=>run);

	-- d987d
	sted987d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord987d,
			Enable=>Enabled987d,
			match=>matchd987d,
			run=>run);

	Enabled987d <= matchd987d OR matchd986d;
	-- d988d
	sted988d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord988d,
			Enable=>Enabled988d,
			match=>matchd988d,
			run=>run);

	Enabled988d <= matchd987d;
	-- d989d
	sted989d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord989d,
			Enable=>Enabled989d,
			match=>matchd989d,
			run=>run);

	Enabled989d <= matchd988d;
	-- d990d
	sted990d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord990d,
			Enable=>Enabled990d,
			match=>matchd990d,
			run=>run);

	Enabled990d <= matchd989d;
	-- d991d
	sted991d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord991d,
			Enable=>Enabled991d,
			match=>matchd991d,
			run=>run);

	Enabled991d <= matchd990d;
	-- d992d
	sted992d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord992d,
			Enable=>Enabled992d,
			match=>matchd992d,
			run=>run);

	Enabled992d <= matchd991d;
	-- d993d
	sted993d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord993d,
			Enable=>Enabled993d,
			match=>matchd993d,
			run=>run);

	Enabled993d <= matchd992d;
	-- d994d
	sted994d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord994d,
			Enable=>Enabled994d,
			match=>matchd994d,
			run=>run);

	Enabled994d <= matchd993d;
	-- d995d
	sted995d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord995d,
			Enable=>Enabled995d,
			match=>matchd995d,
			run=>run);

	Enabled995d <= matchd994d;
	-- d996d
	sted996d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord996d,
			Enable=>Enabled996d,
			match=>matchd996d,
			run=>run);

	Enabled996d <= matchd996d OR matchd995d;
	-- d997d
	sted997d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord997d,
			Enable=>Enabled997d,
			match=>matchd997d,
			run=>run);

	Enabled997d <= matchd996d;
	-- d998d
	sted998d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord998d,
			Enable=>Enabled998d,
			match=>matchd998d,
			run=>run);

	Enabled998d <= matchd997d;
	-- d999d
	sted999d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord999d,
			Enable=>Enabled999d,
			match=>matchd999d,
			run=>run);

	Enabled999d <= matchd998d;
	-- d1000d
	sted1000d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1000d,
			Enable=>Enabled1000d,
			match=>matchd1000d,
			run=>run);

	Enabled1000d <= matchd999d;
	-- d1001d
	sted1001d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1001d,
			Enable=>Enabled1001d,
			match=>matchd1001d,
			run=>run);

	Enabled1001d <= matchd1000d;
	-- d1002d
	sted1002d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1002d,
			Enable=>Enabled1002d,
			match=>matchd1002d,
			run=>run);

	Enabled1002d <= matchd1002d OR matchd1001d;
	-- d1003d
	sted1003d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1003d,
			Enable=>Enabled1003d,
			match=>matchd1003d,
			run=>run);

	Enabled1003d <= matchd1002d;
	-- d1004d
	sted1004d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1004d,
			Enable=>Enabled1004d,
			match=>matchd1004d,
			run=>run);

	Enabled1004d <= matchd1003d;
	-- d1005d
	sted1005d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1005d,
			Enable=>Enabled1005d,
			match=>matchd1005d,
			run=>run);

	Enabled1005d <= matchd1004d;
	-- d1006d
	sted1006d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1006d,
			Enable=>Enabled1006d,
			match=>matchd1006d,
			run=>run);

	Enabled1006d <= matchd1005d;
	-- d1007d
	sted1007d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1007d,
			Enable=>Enabled1007d,
			match=>matchd1007d,
			run=>run);

	reports(40) <= matchd1007d;
	Enabled1007d <= matchd1006d;
	-- d1008d
	sted1008d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1008d,
			Enable=>Enabled1008d,
			match=>matchd1008d,
			run=>run);

	-- d1009d
	sted1009d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1009d,
			Enable=>Enabled1009d,
			match=>matchd1009d,
			run=>run);

	Enabled1009d <= matchd1008d OR matchd1009d;
	-- d1010d
	sted1010d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1010d,
			Enable=>Enabled1010d,
			match=>matchd1010d,
			run=>run);

	Enabled1010d <= matchd1009d;
	-- d1011d
	sted1011d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1011d,
			Enable=>Enabled1011d,
			match=>matchd1011d,
			run=>run);

	Enabled1011d <= matchd1010d;
	-- d1012d
	sted1012d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1012d,
			Enable=>Enabled1012d,
			match=>matchd1012d,
			run=>run);

	Enabled1012d <= matchd1011d;
	-- d1013d
	sted1013d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1013d,
			Enable=>Enabled1013d,
			match=>matchd1013d,
			run=>run);

	Enabled1013d <= matchd1012d;
	-- d1014d
	sted1014d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1014d,
			Enable=>Enabled1014d,
			match=>matchd1014d,
			run=>run);

	Enabled1014d <= matchd1013d;
	-- d1015d
	sted1015d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1015d,
			Enable=>Enabled1015d,
			match=>matchd1015d,
			run=>run);

	Enabled1015d <= matchd1014d;
	-- d1016d
	sted1016d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1016d,
			Enable=>Enabled1016d,
			match=>matchd1016d,
			run=>run);

	Enabled1016d <= matchd1015d;
	-- d1017d
	sted1017d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1017d,
			Enable=>Enabled1017d,
			match=>matchd1017d,
			run=>run);

	Enabled1017d <= matchd1016d;
	-- d1018d
	sted1018d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1018d,
			Enable=>Enabled1018d,
			match=>matchd1018d,
			run=>run);

	Enabled1018d <= matchd1017d OR matchd1018d;
	-- d1019d
	sted1019d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1019d,
			Enable=>Enabled1019d,
			match=>matchd1019d,
			run=>run);

	Enabled1019d <= matchd1018d;
	-- d1020d
	sted1020d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1020d,
			Enable=>Enabled1020d,
			match=>matchd1020d,
			run=>run);

	Enabled1020d <= matchd1019d;
	-- d1021d
	sted1021d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1021d,
			Enable=>Enabled1021d,
			match=>matchd1021d,
			run=>run);

	Enabled1021d <= matchd1020d;
	-- d1022d
	sted1022d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1022d,
			Enable=>Enabled1022d,
			match=>matchd1022d,
			run=>run);

	Enabled1022d <= matchd1021d;
	-- d1023d
	sted1023d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1023d,
			Enable=>Enabled1023d,
			match=>matchd1023d,
			run=>run);

	Enabled1023d <= matchd1022d;
	-- d1024d
	sted1024d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1024d,
			Enable=>Enabled1024d,
			match=>matchd1024d,
			run=>run);

	Enabled1024d <= matchd1024d OR matchd1023d;
	-- d1025d
	sted1025d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1025d,
			Enable=>Enabled1025d,
			match=>matchd1025d,
			run=>run);

	Enabled1025d <= matchd1024d;
	-- d1026d
	sted1026d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1026d,
			Enable=>Enabled1026d,
			match=>matchd1026d,
			run=>run);

	Enabled1026d <= matchd1025d;
	-- d1027d
	sted1027d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1027d,
			Enable=>Enabled1027d,
			match=>matchd1027d,
			run=>run);

	Enabled1027d <= matchd1026d;
	-- d1028d
	sted1028d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1028d,
			Enable=>Enabled1028d,
			match=>matchd1028d,
			run=>run);

	reports(41) <= matchd1028d;
	Enabled1028d <= matchd1027d;
	-- d1029d
	sted1029d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1029d,
			Enable=>Enabled1029d,
			match=>matchd1029d,
			run=>run);

	-- d1030d
	sted1030d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1030d,
			Enable=>Enabled1030d,
			match=>matchd1030d,
			run=>run);

	Enabled1030d <= matchd1029d OR matchd1030d;
	-- d1031d
	sted1031d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1031d,
			Enable=>Enabled1031d,
			match=>matchd1031d,
			run=>run);

	Enabled1031d <= matchd1030d;
	-- d1032d
	sted1032d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1032d,
			Enable=>Enabled1032d,
			match=>matchd1032d,
			run=>run);

	Enabled1032d <= matchd1031d;
	-- d1033d
	sted1033d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1033d,
			Enable=>Enabled1033d,
			match=>matchd1033d,
			run=>run);

	Enabled1033d <= matchd1032d;
	-- d1034d
	sted1034d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1034d,
			Enable=>Enabled1034d,
			match=>matchd1034d,
			run=>run);

	Enabled1034d <= matchd1033d;
	-- d1035d
	sted1035d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1035d,
			Enable=>Enabled1035d,
			match=>matchd1035d,
			run=>run);

	Enabled1035d <= matchd1034d OR matchd1035d;
	-- d1036d
	sted1036d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1036d,
			Enable=>Enabled1036d,
			match=>matchd1036d,
			run=>run);

	Enabled1036d <= matchd1035d;
	-- d1037d
	sted1037d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1037d,
			Enable=>Enabled1037d,
			match=>matchd1037d,
			run=>run);

	Enabled1037d <= matchd1036d;
	-- d1038d
	sted1038d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1038d,
			Enable=>Enabled1038d,
			match=>matchd1038d,
			run=>run);

	Enabled1038d <= matchd1037d;
	-- d1039d
	sted1039d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1039d,
			Enable=>Enabled1039d,
			match=>matchd1039d,
			run=>run);

	reports(42) <= matchd1039d;
	Enabled1039d <= matchd1038d;
	-- d1040d
	sted1040d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1040d,
			Enable=>Enabled1040d,
			match=>matchd1040d,
			run=>run);

	-- d1041d
	sted1041d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1041d,
			Enable=>Enabled1041d,
			match=>matchd1041d,
			run=>run);

	Enabled1041d <= matchd1041d OR matchd1040d;
	-- d1042d
	sted1042d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1042d,
			Enable=>Enabled1042d,
			match=>matchd1042d,
			run=>run);

	Enabled1042d <= matchd1041d;
	-- d1043d
	sted1043d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1043d,
			Enable=>Enabled1043d,
			match=>matchd1043d,
			run=>run);

	Enabled1043d <= matchd1042d;
	-- d1044d
	sted1044d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1044d,
			Enable=>Enabled1044d,
			match=>matchd1044d,
			run=>run);

	Enabled1044d <= matchd1043d;
	-- d1045d
	sted1045d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1045d,
			Enable=>Enabled1045d,
			match=>matchd1045d,
			run=>run);

	Enabled1045d <= matchd1044d;
	-- d1046d
	sted1046d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1046d,
			Enable=>Enabled1046d,
			match=>matchd1046d,
			run=>run);

	Enabled1046d <= matchd1046d OR matchd1045d;
	-- d1047d
	sted1047d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1047d,
			Enable=>Enabled1047d,
			match=>matchd1047d,
			run=>run);

	Enabled1047d <= matchd1046d;
	-- d1048d
	sted1048d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1048d,
			Enable=>Enabled1048d,
			match=>matchd1048d,
			run=>run);

	Enabled1048d <= matchd1047d;
	-- d1049d
	sted1049d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1049d,
			Enable=>Enabled1049d,
			match=>matchd1049d,
			run=>run);

	Enabled1049d <= matchd1048d;
	-- d1050d
	sted1050d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1050d,
			Enable=>Enabled1050d,
			match=>matchd1050d,
			run=>run);

	Enabled1050d <= matchd1049d;
	-- d1051d
	sted1051d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1051d,
			Enable=>Enabled1051d,
			match=>matchd1051d,
			run=>run);

	reports(43) <= matchd1051d;
	Enabled1051d <= matchd1050d;
	-- d1052d
	sted1052d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1052d,
			Enable=>Enabled1052d,
			match=>matchd1052d,
			run=>run);

	-- d1053d
	sted1053d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1053d,
			Enable=>Enabled1053d,
			match=>matchd1053d,
			run=>run);

	Enabled1053d <= matchd1052d OR matchd1053d;
	-- d1054d
	sted1054d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1054d,
			Enable=>Enabled1054d,
			match=>matchd1054d,
			run=>run);

	Enabled1054d <= matchd1053d;
	-- d1055d
	sted1055d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1055d,
			Enable=>Enabled1055d,
			match=>matchd1055d,
			run=>run);

	Enabled1055d <= matchd1054d;
	-- d1056d
	sted1056d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1056d,
			Enable=>Enabled1056d,
			match=>matchd1056d,
			run=>run);

	Enabled1056d <= matchd1055d;
	-- d1057d
	sted1057d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1057d,
			Enable=>Enabled1057d,
			match=>matchd1057d,
			run=>run);

	Enabled1057d <= matchd1056d;
	-- d1058d
	sted1058d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1058d,
			Enable=>Enabled1058d,
			match=>matchd1058d,
			run=>run);

	Enabled1058d <= matchd1057d;
	-- d1059d
	sted1059d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1059d,
			Enable=>Enabled1059d,
			match=>matchd1059d,
			run=>run);

	Enabled1059d <= matchd1058d OR matchd1059d;
	-- d1060d
	sted1060d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1060d,
			Enable=>Enabled1060d,
			match=>matchd1060d,
			run=>run);

	Enabled1060d <= matchd1059d;
	-- d1061d
	sted1061d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1061d,
			Enable=>Enabled1061d,
			match=>matchd1061d,
			run=>run);

	Enabled1061d <= matchd1060d;
	-- d1062d
	sted1062d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1062d,
			Enable=>Enabled1062d,
			match=>matchd1062d,
			run=>run);

	Enabled1062d <= matchd1061d;
	-- d1063d
	sted1063d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1063d,
			Enable=>Enabled1063d,
			match=>matchd1063d,
			run=>run);

	reports(44) <= matchd1063d;
	Enabled1063d <= matchd1062d;
	-- d1064d
	sted1064d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1064d,
			Enable=>Enabled1064d,
			match=>matchd1064d,
			run=>run);

	-- d1065d
	sted1065d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1065d,
			Enable=>Enabled1065d,
			match=>matchd1065d,
			run=>run);

	Enabled1065d <= matchd1065d OR matchd1064d;
	-- d1066d
	sted1066d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1066d,
			Enable=>Enabled1066d,
			match=>matchd1066d,
			run=>run);

	Enabled1066d <= matchd1065d;
	-- d1067d
	sted1067d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1067d,
			Enable=>Enabled1067d,
			match=>matchd1067d,
			run=>run);

	Enabled1067d <= matchd1066d;
	-- d1068d
	sted1068d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1068d,
			Enable=>Enabled1068d,
			match=>matchd1068d,
			run=>run);

	Enabled1068d <= matchd1067d;
	-- d1069d
	sted1069d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1069d,
			Enable=>Enabled1069d,
			match=>matchd1069d,
			run=>run);

	Enabled1069d <= matchd1068d;
	-- d1070d
	sted1070d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1070d,
			Enable=>Enabled1070d,
			match=>matchd1070d,
			run=>run);

	Enabled1070d <= matchd1070d OR matchd1069d;
	-- d1071d
	sted1071d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1071d,
			Enable=>Enabled1071d,
			match=>matchd1071d,
			run=>run);

	Enabled1071d <= matchd1070d;
	-- d1072d
	sted1072d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1072d,
			Enable=>Enabled1072d,
			match=>matchd1072d,
			run=>run);

	Enabled1072d <= matchd1071d;
	-- d1073d
	sted1073d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1073d,
			Enable=>Enabled1073d,
			match=>matchd1073d,
			run=>run);

	Enabled1073d <= matchd1072d;
	-- d1074d
	sted1074d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1074d,
			Enable=>Enabled1074d,
			match=>matchd1074d,
			run=>run);

	Enabled1074d <= matchd1073d;
	-- d1075d
	sted1075d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1075d,
			Enable=>Enabled1075d,
			match=>matchd1075d,
			run=>run);

	reports(45) <= matchd1075d;
	Enabled1075d <= matchd1074d;
	-- d1076d
	sted1076d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1076d,
			Enable=>Enabled1076d,
			match=>matchd1076d,
			run=>run);

	-- d1077d
	sted1077d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1077d,
			Enable=>Enabled1077d,
			match=>matchd1077d,
			run=>run);

	Enabled1077d <= matchd1076d;
	-- d1078d
	sted1078d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1078d,
			Enable=>Enabled1078d,
			match=>matchd1078d,
			run=>run);

	Enabled1078d <= matchd1077d;
	-- d1079d
	sted1079d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1079d,
			Enable=>Enabled1079d,
			match=>matchd1079d,
			run=>run);

	Enabled1079d <= matchd1078d;
	-- d1080d
	sted1080d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1080d,
			Enable=>Enabled1080d,
			match=>matchd1080d,
			run=>run);

	Enabled1080d <= matchd1079d;
	-- d1081d
	sted1081d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1081d,
			Enable=>Enabled1081d,
			match=>matchd1081d,
			run=>run);

	Enabled1081d <= matchd1080d;
	-- d1082d
	sted1082d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1082d,
			Enable=>Enabled1082d,
			match=>matchd1082d,
			run=>run);

	Enabled1082d <= matchd1081d;
	-- d1083d
	sted1083d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1083d,
			Enable=>Enabled1083d,
			match=>matchd1083d,
			run=>run);

	Enabled1083d <= matchd1082d;
	-- d1084d
	sted1084d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1084d,
			Enable=>Enabled1084d,
			match=>matchd1084d,
			run=>run);

	reports(46) <= matchd1084d;
	Enabled1084d <= matchd1083d;
	-- d1085d
	sted1085d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1085d,
			Enable=>Enabled1085d,
			match=>matchd1085d,
			run=>run);

	-- d1086d
	sted1086d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1086d,
			Enable=>Enabled1086d,
			match=>matchd1086d,
			run=>run);

	Enabled1086d <= matchd1086d OR matchd1085d;
	-- d1087d
	sted1087d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1087d,
			Enable=>Enabled1087d,
			match=>matchd1087d,
			run=>run);

	Enabled1087d <= matchd1086d;
	-- d1088d
	sted1088d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1088d,
			Enable=>Enabled1088d,
			match=>matchd1088d,
			run=>run);

	Enabled1088d <= matchd1087d OR matchd1088d;
	-- d1089d
	sted1089d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1089d,
			Enable=>Enabled1089d,
			match=>matchd1089d,
			run=>run);

	Enabled1089d <= matchd1088d;
	-- d1090d
	sted1090d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1090d,
			Enable=>Enabled1090d,
			match=>matchd1090d,
			run=>run);

	Enabled1090d <= matchd1090d OR matchd1089d;
	-- d1091d
	sted1091d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1091d,
			Enable=>Enabled1091d,
			match=>matchd1091d,
			run=>run);

	Enabled1091d <= matchd1090d;
	-- d1092d
	sted1092d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1092d,
			Enable=>Enabled1092d,
			match=>matchd1092d,
			run=>run);

	Enabled1092d <= matchd1091d;
	-- d1093d
	sted1093d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1093d,
			Enable=>Enabled1093d,
			match=>matchd1093d,
			run=>run);

	Enabled1093d <= matchd1092d;
	-- d1094d
	sted1094d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1094d,
			Enable=>Enabled1094d,
			match=>matchd1094d,
			run=>run);

	Enabled1094d <= matchd1093d;
	-- d1095d
	sted1095d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1095d,
			Enable=>Enabled1095d,
			match=>matchd1095d,
			run=>run);

	Enabled1095d <= matchd1094d;
	-- d1096d
	sted1096d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1096d,
			Enable=>Enabled1096d,
			match=>matchd1096d,
			run=>run);

	Enabled1096d <= matchd1095d OR matchd1096d;
	-- d1097d
	sted1097d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1097d,
			Enable=>Enabled1097d,
			match=>matchd1097d,
			run=>run);

	Enabled1097d <= matchd1096d;
	-- d1098d
	sted1098d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1098d,
			Enable=>Enabled1098d,
			match=>matchd1098d,
			run=>run);

	Enabled1098d <= matchd1097d;
	-- d1099d
	sted1099d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1099d,
			Enable=>Enabled1099d,
			match=>matchd1099d,
			run=>run);

	Enabled1099d <= matchd1098d;
	-- d1100d
	sted1100d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1100d,
			Enable=>Enabled1100d,
			match=>matchd1100d,
			run=>run);

	Enabled1100d <= matchd1099d;
	-- d1101d
	sted1101d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1101d,
			Enable=>Enabled1101d,
			match=>matchd1101d,
			run=>run);

	Enabled1101d <= matchd1100d;
	-- d1102d
	sted1102d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1102d,
			Enable=>Enabled1102d,
			match=>matchd1102d,
			run=>run);

	-- d1103d
	sted1103d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1103d,
			Enable=>Enabled1103d,
			match=>matchd1103d,
			run=>run);

	Enabled1103d <= matchd1102d OR matchd1103d;
	-- d1104d
	sted1104d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1104d,
			Enable=>Enabled1104d,
			match=>matchd1104d,
			run=>run);

	Enabled1104d <= matchd1103d;
	-- d1105d
	sted1105d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1105d,
			Enable=>Enabled1105d,
			match=>matchd1105d,
			run=>run);

	Enabled1105d <= matchd1104d;
	-- d1106d
	sted1106d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1106d,
			Enable=>Enabled1106d,
			match=>matchd1106d,
			run=>run);

	Enabled1106d <= matchd1105d;
	-- d1107d
	sted1107d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1107d,
			Enable=>Enabled1107d,
			match=>matchd1107d,
			run=>run);

	Enabled1107d <= matchd1106d;
	-- d1108d
	sted1108d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1108d,
			Enable=>Enabled1108d,
			match=>matchd1108d,
			run=>run);

	Enabled1108d <= matchd1107d;
	-- d1109d
	sted1109d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1109d,
			Enable=>Enabled1109d,
			match=>matchd1109d,
			run=>run);

	Enabled1109d <= matchd1108d OR matchd1109d;
	-- d1110d
	sted1110d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1110d,
			Enable=>Enabled1110d,
			match=>matchd1110d,
			run=>run);

	Enabled1110d <= matchd1109d;
	-- d1111d
	sted1111d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1111d,
			Enable=>Enabled1111d,
			match=>matchd1111d,
			run=>run);

	Enabled1111d <= matchd1111d OR matchd1110d;
	-- d1112d
	sted1112d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1112d,
			Enable=>Enabled1112d,
			match=>matchd1112d,
			run=>run);

	Enabled1112d <= matchd1111d;
	-- d1113d
	sted1113d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1113d,
			Enable=>Enabled1113d,
			match=>matchd1113d,
			run=>run);

	Enabled1113d <= matchd1113d OR matchd1112d;
	-- d1114d
	sted1114d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1114d,
			Enable=>Enabled1114d,
			match=>matchd1114d,
			run=>run);

	Enabled1114d <= matchd1113d;
	-- d1115d
	sted1115d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1115d,
			Enable=>Enabled1115d,
			match=>matchd1115d,
			run=>run);

	Enabled1115d <= matchd1114d;
	-- d1116d
	sted1116d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1116d,
			Enable=>Enabled1116d,
			match=>matchd1116d,
			run=>run);

	Enabled1116d <= matchd1115d;
	-- d1117d
	sted1117d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1117d,
			Enable=>Enabled1117d,
			match=>matchd1117d,
			run=>run);

	Enabled1117d <= matchd1116d;
	-- d1118d
	sted1118d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1118d,
			Enable=>Enabled1118d,
			match=>matchd1118d,
			run=>run);

	Enabled1118d <= matchd1117d;
	-- d1120d
	sted1120d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1120d,
			Enable=>Enabled1120d,
			match=>matchd1120d,
			run=>run);

	-- d1121d
	sted1121d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1121d,
			Enable=>Enabled1121d,
			match=>matchd1121d,
			run=>run);

	Enabled1121d <= matchd1120d OR matchd1121d;
	-- d1122d
	sted1122d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1122d,
			Enable=>Enabled1122d,
			match=>matchd1122d,
			run=>run);

	Enabled1122d <= matchd1121d;
	-- d1123d
	sted1123d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1123d,
			Enable=>Enabled1123d,
			match=>matchd1123d,
			run=>run);

	Enabled1123d <= matchd1122d;
	-- d1124d
	sted1124d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1124d,
			Enable=>Enabled1124d,
			match=>matchd1124d,
			run=>run);

	Enabled1124d <= matchd1123d;
	-- d1125d
	sted1125d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1125d,
			Enable=>Enabled1125d,
			match=>matchd1125d,
			run=>run);

	Enabled1125d <= matchd1124d;
	-- d1126d
	sted1126d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1126d,
			Enable=>Enabled1126d,
			match=>matchd1126d,
			run=>run);

	Enabled1126d <= matchd1125d OR matchd1126d;
	-- d1127d
	sted1127d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1127d,
			Enable=>Enabled1127d,
			match=>matchd1127d,
			run=>run);

	Enabled1127d <= matchd1126d;
	-- d1128d
	sted1128d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1128d,
			Enable=>Enabled1128d,
			match=>matchd1128d,
			run=>run);

	Enabled1128d <= matchd1127d;
	-- d1129d
	sted1129d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1129d,
			Enable=>Enabled1129d,
			match=>matchd1129d,
			run=>run);

	Enabled1129d <= matchd1128d;
	-- d1130d
	sted1130d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1130d,
			Enable=>Enabled1130d,
			match=>matchd1130d,
			run=>run);

	reports(47) <= matchd1130d;
	Enabled1130d <= matchd1129d;
	-- d1131d
	sted1131d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1131d,
			Enable=>Enabled1131d,
			match=>matchd1131d,
			run=>run);

	-- d1132d
	sted1132d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1132d,
			Enable=>Enabled1132d,
			match=>matchd1132d,
			run=>run);

	Enabled1132d <= matchd1131d OR matchd1132d;
	-- d1133d
	sted1133d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1133d,
			Enable=>Enabled1133d,
			match=>matchd1133d,
			run=>run);

	Enabled1133d <= matchd1132d;
	-- d1134d
	sted1134d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1134d,
			Enable=>Enabled1134d,
			match=>matchd1134d,
			run=>run);

	Enabled1134d <= matchd1133d;
	-- d1135d
	sted1135d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1135d,
			Enable=>Enabled1135d,
			match=>matchd1135d,
			run=>run);

	Enabled1135d <= matchd1134d;
	-- d1136d
	sted1136d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1136d,
			Enable=>Enabled1136d,
			match=>matchd1136d,
			run=>run);

	Enabled1136d <= matchd1135d;
	-- d1137d
	sted1137d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1137d,
			Enable=>Enabled1137d,
			match=>matchd1137d,
			run=>run);

	Enabled1137d <= matchd1136d;
	-- d1138d
	sted1138d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1138d,
			Enable=>Enabled1138d,
			match=>matchd1138d,
			run=>run);

	Enabled1138d <= matchd1138d OR matchd1137d;
	-- d1139d
	sted1139d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1139d,
			Enable=>Enabled1139d,
			match=>matchd1139d,
			run=>run);

	Enabled1139d <= matchd1138d;
	-- d1140d
	sted1140d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1140d,
			Enable=>Enabled1140d,
			match=>matchd1140d,
			run=>run);

	Enabled1140d <= matchd1139d;
	-- d1141d
	sted1141d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1141d,
			Enable=>Enabled1141d,
			match=>matchd1141d,
			run=>run);

	Enabled1141d <= matchd1140d;
	-- d1142d
	sted1142d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1142d,
			Enable=>Enabled1142d,
			match=>matchd1142d,
			run=>run);

	reports(48) <= matchd1142d;
	Enabled1142d <= matchd1141d;
	-- d1143d
	sted1143d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1143d,
			Enable=>Enabled1143d,
			match=>matchd1143d,
			run=>run);

	-- d1144d
	sted1144d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1144d,
			Enable=>Enabled1144d,
			match=>matchd1144d,
			run=>run);

	Enabled1144d <= matchd1143d;
	-- d1145d
	sted1145d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1145d,
			Enable=>Enabled1145d,
			match=>matchd1145d,
			run=>run);

	Enabled1145d <= matchd1144d;
	-- d1146d
	sted1146d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1146d,
			Enable=>Enabled1146d,
			match=>matchd1146d,
			run=>run);

	Enabled1146d <= matchd1145d;
	-- d1147d
	sted1147d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1147d,
			Enable=>Enabled1147d,
			match=>matchd1147d,
			run=>run);

	Enabled1147d <= matchd1146d;
	-- d1148d
	sted1148d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1148d,
			Enable=>Enabled1148d,
			match=>matchd1148d,
			run=>run);

	Enabled1148d <= matchd1147d;
	-- d1149d
	sted1149d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1149d,
			Enable=>Enabled1149d,
			match=>matchd1149d,
			run=>run);

	Enabled1149d <= matchd1148d;
	-- d1150d
	sted1150d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1150d,
			Enable=>Enabled1150d,
			match=>matchd1150d,
			run=>run);

	Enabled1150d <= matchd1149d;
	-- d1151d
	sted1151d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1151d,
			Enable=>Enabled1151d,
			match=>matchd1151d,
			run=>run);

	Enabled1151d <= matchd1150d;
	-- d1152d
	sted1152d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1152d,
			Enable=>Enabled1152d,
			match=>matchd1152d,
			run=>run);

	reports(49) <= matchd1152d;
	Enabled1152d <= matchd1151d;
	-- d1153d
	sted1153d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1153d,
			Enable=>Enabled1153d,
			match=>matchd1153d,
			run=>run);

	-- d1154d
	sted1154d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1154d,
			Enable=>Enabled1154d,
			match=>matchd1154d,
			run=>run);

	Enabled1154d <= matchd1153d OR matchd1154d;
	-- d1155d
	sted1155d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1155d,
			Enable=>Enabled1155d,
			match=>matchd1155d,
			run=>run);

	Enabled1155d <= matchd1154d;
	-- d1156d
	sted1156d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1156d,
			Enable=>Enabled1156d,
			match=>matchd1156d,
			run=>run);

	Enabled1156d <= matchd1155d;
	-- d1157d
	sted1157d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1157d,
			Enable=>Enabled1157d,
			match=>matchd1157d,
			run=>run);

	Enabled1157d <= matchd1156d;
	-- d1158d
	sted1158d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1158d,
			Enable=>Enabled1158d,
			match=>matchd1158d,
			run=>run);

	Enabled1158d <= matchd1157d;
	-- d1159d
	sted1159d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1159d,
			Enable=>Enabled1159d,
			match=>matchd1159d,
			run=>run);

	Enabled1159d <= matchd1159d OR matchd1158d;
	-- d1160d
	sted1160d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1160d,
			Enable=>Enabled1160d,
			match=>matchd1160d,
			run=>run);

	Enabled1160d <= matchd1159d;
	-- d1161d
	sted1161d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1161d,
			Enable=>Enabled1161d,
			match=>matchd1161d,
			run=>run);

	Enabled1161d <= matchd1160d OR matchd1161d;
	-- d1162d
	sted1162d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1162d,
			Enable=>Enabled1162d,
			match=>matchd1162d,
			run=>run);

	Enabled1162d <= matchd1161d;
	-- d1163d
	sted1163d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1163d,
			Enable=>Enabled1163d,
			match=>matchd1163d,
			run=>run);

	Enabled1163d <= matchd1162d OR matchd1163d;
	-- d1164d
	sted1164d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1164d,
			Enable=>Enabled1164d,
			match=>matchd1164d,
			run=>run);

	Enabled1164d <= matchd1163d;
	-- d1165d
	sted1165d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1165d,
			Enable=>Enabled1165d,
			match=>matchd1165d,
			run=>run);

	Enabled1165d <= matchd1164d;
	-- d1166d
	sted1166d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1166d,
			Enable=>Enabled1166d,
			match=>matchd1166d,
			run=>run);

	Enabled1166d <= matchd1165d;
	-- d1167d
	sted1167d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1167d,
			Enable=>Enabled1167d,
			match=>matchd1167d,
			run=>run);

	Enabled1167d <= matchd1166d;
	-- d1168d
	sted1168d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1168d,
			Enable=>Enabled1168d,
			match=>matchd1168d,
			run=>run);

	reports(50) <= matchd1168d;
	Enabled1168d <= matchd1167d;
	-- d1169d
	sted1169d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1169d,
			Enable=>Enabled1169d,
			match=>matchd1169d,
			run=>run);

	-- d1170d
	sted1170d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1170d,
			Enable=>Enabled1170d,
			match=>matchd1170d,
			run=>run);

	Enabled1170d <= matchd1169d;
	-- d1171d
	sted1171d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1171d,
			Enable=>Enabled1171d,
			match=>matchd1171d,
			run=>run);

	Enabled1171d <= matchd1170d;
	-- d1172d
	sted1172d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1172d,
			Enable=>Enabled1172d,
			match=>matchd1172d,
			run=>run);

	Enabled1172d <= matchd1171d;
	-- d1173d
	sted1173d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1173d,
			Enable=>Enabled1173d,
			match=>matchd1173d,
			run=>run);

	Enabled1173d <= matchd1172d;
	-- d1174d
	sted1174d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1174d,
			Enable=>Enabled1174d,
			match=>matchd1174d,
			run=>run);

	Enabled1174d <= matchd1173d;
	-- d1175d
	sted1175d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1175d,
			Enable=>Enabled1175d,
			match=>matchd1175d,
			run=>run);

	Enabled1175d <= matchd1174d;
	-- d1176d
	sted1176d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1176d,
			Enable=>Enabled1176d,
			match=>matchd1176d,
			run=>run);

	Enabled1176d <= matchd1176d OR matchd1175d;
	-- d1177d
	sted1177d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1177d,
			Enable=>Enabled1177d,
			match=>matchd1177d,
			run=>run);

	Enabled1177d <= matchd1176d;
	-- d1178d
	sted1178d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1178d,
			Enable=>Enabled1178d,
			match=>matchd1178d,
			run=>run);

	Enabled1178d <= matchd1177d;
	-- d1179d
	sted1179d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1179d,
			Enable=>Enabled1179d,
			match=>matchd1179d,
			run=>run);

	Enabled1179d <= matchd1178d;
	-- d1180d
	sted1180d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1180d,
			Enable=>Enabled1180d,
			match=>matchd1180d,
			run=>run);

	Enabled1180d <= matchd1179d;
	-- d1181d
	sted1181d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1181d,
			Enable=>Enabled1181d,
			match=>matchd1181d,
			run=>run);

	reports(51) <= matchd1181d;
	Enabled1181d <= matchd1180d;
	-- d1182d
	sted1182d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1182d,
			Enable=>Enabled1182d,
			match=>matchd1182d,
			run=>run);

	-- d1183d
	sted1183d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1183d,
			Enable=>Enabled1183d,
			match=>matchd1183d,
			run=>run);

	Enabled1183d <= matchd1182d OR matchd1183d;
	-- d1184d
	sted1184d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1184d,
			Enable=>Enabled1184d,
			match=>matchd1184d,
			run=>run);

	Enabled1184d <= matchd1183d;
	-- d1185d
	sted1185d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1185d,
			Enable=>Enabled1185d,
			match=>matchd1185d,
			run=>run);

	Enabled1185d <= matchd1184d;
	-- d1186d
	sted1186d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1186d,
			Enable=>Enabled1186d,
			match=>matchd1186d,
			run=>run);

	Enabled1186d <= matchd1185d;
	-- d1187d
	sted1187d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1187d,
			Enable=>Enabled1187d,
			match=>matchd1187d,
			run=>run);

	Enabled1187d <= matchd1186d;
	-- d1188d
	sted1188d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1188d,
			Enable=>Enabled1188d,
			match=>matchd1188d,
			run=>run);

	Enabled1188d <= matchd1188d OR matchd1187d;
	-- d1189d
	sted1189d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1189d,
			Enable=>Enabled1189d,
			match=>matchd1189d,
			run=>run);

	Enabled1189d <= matchd1188d;
	-- d1190d
	sted1190d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1190d,
			Enable=>Enabled1190d,
			match=>matchd1190d,
			run=>run);

	Enabled1190d <= matchd1189d;
	-- d1191d
	sted1191d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1191d,
			Enable=>Enabled1191d,
			match=>matchd1191d,
			run=>run);

	Enabled1191d <= matchd1190d;
	-- d1192d
	sted1192d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1192d,
			Enable=>Enabled1192d,
			match=>matchd1192d,
			run=>run);

	reports(52) <= matchd1192d;
	Enabled1192d <= matchd1191d;
	-- d1193d
	sted1193d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1193d,
			Enable=>Enabled1193d,
			match=>matchd1193d,
			run=>run);

	-- d1194d
	sted1194d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1194d,
			Enable=>Enabled1194d,
			match=>matchd1194d,
			run=>run);

	Enabled1194d <= matchd1193d OR matchd1194d;
	-- d1195d
	sted1195d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1195d,
			Enable=>Enabled1195d,
			match=>matchd1195d,
			run=>run);

	Enabled1195d <= matchd1194d;
	-- d1196d
	sted1196d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1196d,
			Enable=>Enabled1196d,
			match=>matchd1196d,
			run=>run);

	Enabled1196d <= matchd1195d;
	-- d1197d
	sted1197d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1197d,
			Enable=>Enabled1197d,
			match=>matchd1197d,
			run=>run);

	Enabled1197d <= matchd1196d;
	-- d1198d
	sted1198d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1198d,
			Enable=>Enabled1198d,
			match=>matchd1198d,
			run=>run);

	Enabled1198d <= matchd1197d;
	-- d1199d
	sted1199d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1199d,
			Enable=>Enabled1199d,
			match=>matchd1199d,
			run=>run);

	Enabled1199d <= matchd1198d;
	-- d1200d
	sted1200d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1200d,
			Enable=>Enabled1200d,
			match=>matchd1200d,
			run=>run);

	Enabled1200d <= matchd1199d;
	-- d1201d
	sted1201d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1201d,
			Enable=>Enabled1201d,
			match=>matchd1201d,
			run=>run);

	Enabled1201d <= matchd1200d;
	-- d1202d
	sted1202d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1202d,
			Enable=>Enabled1202d,
			match=>matchd1202d,
			run=>run);

	Enabled1202d <= matchd1201d;
	-- d1203d
	sted1203d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1203d,
			Enable=>Enabled1203d,
			match=>matchd1203d,
			run=>run);

	Enabled1203d <= matchd1203d OR matchd1202d;
	-- d1204d
	sted1204d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1204d,
			Enable=>Enabled1204d,
			match=>matchd1204d,
			run=>run);

	Enabled1204d <= matchd1203d;
	-- d1205d
	sted1205d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1205d,
			Enable=>Enabled1205d,
			match=>matchd1205d,
			run=>run);

	Enabled1205d <= matchd1204d;
	-- d1206d
	sted1206d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1206d,
			Enable=>Enabled1206d,
			match=>matchd1206d,
			run=>run);

	Enabled1206d <= matchd1205d;
	-- d1207d
	sted1207d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1207d,
			Enable=>Enabled1207d,
			match=>matchd1207d,
			run=>run);

	Enabled1207d <= matchd1206d;
	-- d1208d
	sted1208d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1208d,
			Enable=>Enabled1208d,
			match=>matchd1208d,
			run=>run);

	Enabled1208d <= matchd1207d;
	-- d1209d
	sted1209d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1209d,
			Enable=>Enabled1209d,
			match=>matchd1209d,
			run=>run);

	Enabled1209d <= matchd1208d OR matchd1209d;
	-- d1210d
	sted1210d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1210d,
			Enable=>Enabled1210d,
			match=>matchd1210d,
			run=>run);

	Enabled1210d <= matchd1209d;
	-- d1211d
	sted1211d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1211d,
			Enable=>Enabled1211d,
			match=>matchd1211d,
			run=>run);

	Enabled1211d <= matchd1210d;
	-- d1212d
	sted1212d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1212d,
			Enable=>Enabled1212d,
			match=>matchd1212d,
			run=>run);

	Enabled1212d <= matchd1211d;
	-- d1213d
	sted1213d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1213d,
			Enable=>Enabled1213d,
			match=>matchd1213d,
			run=>run);

	reports(53) <= matchd1213d;
	Enabled1213d <= matchd1212d;
	-- d1214d
	sted1214d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1214d,
			Enable=>Enabled1214d,
			match=>matchd1214d,
			run=>run);

	-- d1215d
	sted1215d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1215d,
			Enable=>Enabled1215d,
			match=>matchd1215d,
			run=>run);

	Enabled1215d <= matchd1215d OR matchd1214d;
	-- d1216d
	sted1216d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1216d,
			Enable=>Enabled1216d,
			match=>matchd1216d,
			run=>run);

	Enabled1216d <= matchd1215d;
	-- d1217d
	sted1217d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1217d,
			Enable=>Enabled1217d,
			match=>matchd1217d,
			run=>run);

	Enabled1217d <= matchd1216d;
	-- d1218d
	sted1218d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1218d,
			Enable=>Enabled1218d,
			match=>matchd1218d,
			run=>run);

	Enabled1218d <= matchd1217d;
	-- d1219d
	sted1219d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1219d,
			Enable=>Enabled1219d,
			match=>matchd1219d,
			run=>run);

	Enabled1219d <= matchd1218d;
	-- d1220d
	sted1220d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1220d,
			Enable=>Enabled1220d,
			match=>matchd1220d,
			run=>run);

	Enabled1220d <= matchd1219d OR matchd1220d;
	-- d1221d
	sted1221d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1221d,
			Enable=>Enabled1221d,
			match=>matchd1221d,
			run=>run);

	Enabled1221d <= matchd1220d;
	-- d1222d
	sted1222d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1222d,
			Enable=>Enabled1222d,
			match=>matchd1222d,
			run=>run);

	Enabled1222d <= matchd1221d;
	-- d1223d
	sted1223d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1223d,
			Enable=>Enabled1223d,
			match=>matchd1223d,
			run=>run);

	Enabled1223d <= matchd1222d;
	-- d1224d
	sted1224d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1224d,
			Enable=>Enabled1224d,
			match=>matchd1224d,
			run=>run);

	reports(54) <= matchd1224d;
	Enabled1224d <= matchd1223d;
	-- d1225d
	sted1225d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1225d,
			Enable=>Enabled1225d,
			match=>matchd1225d,
			run=>run);

	-- d1226d
	sted1226d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1226d,
			Enable=>Enabled1226d,
			match=>matchd1226d,
			run=>run);

	Enabled1226d <= matchd1226d OR matchd1225d;
	-- d1227d
	sted1227d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1227d,
			Enable=>Enabled1227d,
			match=>matchd1227d,
			run=>run);

	Enabled1227d <= matchd1226d;
	-- d1228d
	sted1228d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1228d,
			Enable=>Enabled1228d,
			match=>matchd1228d,
			run=>run);

	Enabled1228d <= matchd1227d;
	-- d1229d
	sted1229d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1229d,
			Enable=>Enabled1229d,
			match=>matchd1229d,
			run=>run);

	Enabled1229d <= matchd1228d;
	-- d1230d
	sted1230d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1230d,
			Enable=>Enabled1230d,
			match=>matchd1230d,
			run=>run);

	Enabled1230d <= matchd1229d;
	-- d1231d
	sted1231d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1231d,
			Enable=>Enabled1231d,
			match=>matchd1231d,
			run=>run);

	Enabled1231d <= matchd1230d OR matchd1231d;
	-- d1232d
	sted1232d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1232d,
			Enable=>Enabled1232d,
			match=>matchd1232d,
			run=>run);

	Enabled1232d <= matchd1231d;
	-- d1233d
	sted1233d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1233d,
			Enable=>Enabled1233d,
			match=>matchd1233d,
			run=>run);

	Enabled1233d <= matchd1232d;
	-- d1234d
	sted1234d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1234d,
			Enable=>Enabled1234d,
			match=>matchd1234d,
			run=>run);

	Enabled1234d <= matchd1233d;
	-- d1235d
	sted1235d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1235d,
			Enable=>Enabled1235d,
			match=>matchd1235d,
			run=>run);

	Enabled1235d <= matchd1234d;
	-- d1236d
	sted1236d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1236d,
			Enable=>Enabled1236d,
			match=>matchd1236d,
			run=>run);

	Enabled1236d <= matchd1235d;
	-- d1237d
	sted1237d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1237d,
			Enable=>Enabled1237d,
			match=>matchd1237d,
			run=>run);

	Enabled1237d <= matchd1236d OR matchd1237d;
	-- d1238d
	sted1238d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1238d,
			Enable=>Enabled1238d,
			match=>matchd1238d,
			run=>run);

	Enabled1238d <= matchd1237d;
	-- d1239d
	sted1239d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1239d,
			Enable=>Enabled1239d,
			match=>matchd1239d,
			run=>run);

	Enabled1239d <= matchd1238d;
	-- d1240d
	sted1240d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1240d,
			Enable=>Enabled1240d,
			match=>matchd1240d,
			run=>run);

	Enabled1240d <= matchd1239d;
	-- d1241d
	sted1241d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1241d,
			Enable=>Enabled1241d,
			match=>matchd1241d,
			run=>run);

	reports(55) <= matchd1241d;
	Enabled1241d <= matchd1240d;
	-- d1242d
	sted1242d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1242d,
			Enable=>Enabled1242d,
			match=>matchd1242d,
			run=>run);

	-- d1243d
	sted1243d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1243d,
			Enable=>Enabled1243d,
			match=>matchd1243d,
			run=>run);

	Enabled1243d <= matchd1242d OR matchd1243d;
	-- d1244d
	sted1244d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1244d,
			Enable=>Enabled1244d,
			match=>matchd1244d,
			run=>run);

	Enabled1244d <= matchd1243d;
	-- d1245d
	sted1245d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1245d,
			Enable=>Enabled1245d,
			match=>matchd1245d,
			run=>run);

	Enabled1245d <= matchd1244d;
	-- d1246d
	sted1246d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1246d,
			Enable=>Enabled1246d,
			match=>matchd1246d,
			run=>run);

	Enabled1246d <= matchd1245d;
	-- d1247d
	sted1247d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1247d,
			Enable=>Enabled1247d,
			match=>matchd1247d,
			run=>run);

	Enabled1247d <= matchd1246d;
	-- d1248d
	sted1248d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1248d,
			Enable=>Enabled1248d,
			match=>matchd1248d,
			run=>run);

	Enabled1248d <= matchd1247d OR matchd1248d;
	-- d1249d
	sted1249d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1249d,
			Enable=>Enabled1249d,
			match=>matchd1249d,
			run=>run);

	Enabled1249d <= matchd1248d;
	-- d1250d
	sted1250d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1250d,
			Enable=>Enabled1250d,
			match=>matchd1250d,
			run=>run);

	Enabled1250d <= matchd1249d;
	-- d1251d
	sted1251d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1251d,
			Enable=>Enabled1251d,
			match=>matchd1251d,
			run=>run);

	Enabled1251d <= matchd1250d;
	-- d1252d
	sted1252d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1252d,
			Enable=>Enabled1252d,
			match=>matchd1252d,
			run=>run);

	Enabled1252d <= matchd1251d;
	-- d1253d
	sted1253d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1253d,
			Enable=>Enabled1253d,
			match=>matchd1253d,
			run=>run);

	reports(56) <= matchd1253d;
	Enabled1253d <= matchd1252d;
	-- d1254d
	sted1254d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1254d,
			Enable=>Enabled1254d,
			match=>matchd1254d,
			run=>run);

	-- d1255d
	sted1255d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1255d,
			Enable=>Enabled1255d,
			match=>matchd1255d,
			run=>run);

	Enabled1255d <= matchd1255d OR matchd1254d;
	-- d1256d
	sted1256d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1256d,
			Enable=>Enabled1256d,
			match=>matchd1256d,
			run=>run);

	Enabled1256d <= matchd1255d;
	-- d1257d
	sted1257d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1257d,
			Enable=>Enabled1257d,
			match=>matchd1257d,
			run=>run);

	Enabled1257d <= matchd1256d;
	-- d1258d
	sted1258d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1258d,
			Enable=>Enabled1258d,
			match=>matchd1258d,
			run=>run);

	Enabled1258d <= matchd1257d;
	-- d1259d
	sted1259d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1259d,
			Enable=>Enabled1259d,
			match=>matchd1259d,
			run=>run);

	Enabled1259d <= matchd1258d;
	-- d1260d
	sted1260d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1260d,
			Enable=>Enabled1260d,
			match=>matchd1260d,
			run=>run);

	Enabled1260d <= matchd1259d;
	-- d1261d
	sted1261d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1261d,
			Enable=>Enabled1261d,
			match=>matchd1261d,
			run=>run);

	Enabled1261d <= matchd1261d OR matchd1260d;
	-- d1262d
	sted1262d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1262d,
			Enable=>Enabled1262d,
			match=>matchd1262d,
			run=>run);

	Enabled1262d <= matchd1261d;
	-- d1263d
	sted1263d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1263d,
			Enable=>Enabled1263d,
			match=>matchd1263d,
			run=>run);

	Enabled1263d <= matchd1262d;
	-- d1264d
	sted1264d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1264d,
			Enable=>Enabled1264d,
			match=>matchd1264d,
			run=>run);

	Enabled1264d <= matchd1263d;
	-- d1265d
	sted1265d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1265d,
			Enable=>Enabled1265d,
			match=>matchd1265d,
			run=>run);

	Enabled1265d <= matchd1264d;
	-- d1266d
	sted1266d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1266d,
			Enable=>Enabled1266d,
			match=>matchd1266d,
			run=>run);

	reports(57) <= matchd1266d;
	Enabled1266d <= matchd1265d;
	-- d1267d
	sted1267d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1267d,
			Enable=>Enabled1267d,
			match=>matchd1267d,
			run=>run);

	-- d1268d
	sted1268d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1268d,
			Enable=>Enabled1268d,
			match=>matchd1268d,
			run=>run);

	Enabled1268d <= matchd1267d OR matchd1268d;
	-- d1269d
	sted1269d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1269d,
			Enable=>Enabled1269d,
			match=>matchd1269d,
			run=>run);

	Enabled1269d <= matchd1268d;
	-- d1270d
	sted1270d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1270d,
			Enable=>Enabled1270d,
			match=>matchd1270d,
			run=>run);

	Enabled1270d <= matchd1270d OR matchd1269d;
	-- d1271d
	sted1271d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1271d,
			Enable=>Enabled1271d,
			match=>matchd1271d,
			run=>run);

	Enabled1271d <= matchd1270d;
	-- d1272d
	sted1272d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1272d,
			Enable=>Enabled1272d,
			match=>matchd1272d,
			run=>run);

	Enabled1272d <= matchd1271d OR matchd1272d;
	-- d1273d
	sted1273d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1273d,
			Enable=>Enabled1273d,
			match=>matchd1273d,
			run=>run);

	Enabled1273d <= matchd1272d;
	-- d1274d
	sted1274d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1274d,
			Enable=>Enabled1274d,
			match=>matchd1274d,
			run=>run);

	Enabled1274d <= matchd1273d;
	-- d1275d
	sted1275d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1275d,
			Enable=>Enabled1275d,
			match=>matchd1275d,
			run=>run);

	Enabled1275d <= matchd1274d;
	-- d1276d
	sted1276d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1276d,
			Enable=>Enabled1276d,
			match=>matchd1276d,
			run=>run);

	Enabled1276d <= matchd1275d;
	-- d1277d
	sted1277d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1277d,
			Enable=>Enabled1277d,
			match=>matchd1277d,
			run=>run);

	Enabled1277d <= matchd1276d;
	-- d1278d
	sted1278d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1278d,
			Enable=>Enabled1278d,
			match=>matchd1278d,
			run=>run);

	Enabled1278d <= matchd1278d OR matchd1277d;
	-- d1279d
	sted1279d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1279d,
			Enable=>Enabled1279d,
			match=>matchd1279d,
			run=>run);

	Enabled1279d <= matchd1278d;
	-- d1280d
	sted1280d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1280d,
			Enable=>Enabled1280d,
			match=>matchd1280d,
			run=>run);

	Enabled1280d <= matchd1279d;
	-- d1281d
	sted1281d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1281d,
			Enable=>Enabled1281d,
			match=>matchd1281d,
			run=>run);

	Enabled1281d <= matchd1280d;
	-- d1282d
	sted1282d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1282d,
			Enable=>Enabled1282d,
			match=>matchd1282d,
			run=>run);

	Enabled1282d <= matchd1281d;
	-- d1283d
	sted1283d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1283d,
			Enable=>Enabled1283d,
			match=>matchd1283d,
			run=>run);

	-- d1284d
	sted1284d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1284d,
			Enable=>Enabled1284d,
			match=>matchd1284d,
			run=>run);

	Enabled1284d <= matchd1284d OR matchd1283d;
	-- d1285d
	sted1285d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1285d,
			Enable=>Enabled1285d,
			match=>matchd1285d,
			run=>run);

	Enabled1285d <= matchd1284d;
	-- d1286d
	sted1286d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1286d,
			Enable=>Enabled1286d,
			match=>matchd1286d,
			run=>run);

	Enabled1286d <= matchd1285d;
	-- d1287d
	sted1287d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1287d,
			Enable=>Enabled1287d,
			match=>matchd1287d,
			run=>run);

	Enabled1287d <= matchd1286d;
	-- d1288d
	sted1288d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1288d,
			Enable=>Enabled1288d,
			match=>matchd1288d,
			run=>run);

	Enabled1288d <= matchd1287d;
	-- d1289d
	sted1289d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1289d,
			Enable=>Enabled1289d,
			match=>matchd1289d,
			run=>run);

	Enabled1289d <= matchd1288d;
	-- d1290d
	sted1290d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1290d,
			Enable=>Enabled1290d,
			match=>matchd1290d,
			run=>run);

	Enabled1290d <= matchd1290d OR matchd1289d;
	-- d1291d
	sted1291d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1291d,
			Enable=>Enabled1291d,
			match=>matchd1291d,
			run=>run);

	Enabled1291d <= matchd1290d;
	-- d1292d
	sted1292d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1292d,
			Enable=>Enabled1292d,
			match=>matchd1292d,
			run=>run);

	Enabled1292d <= matchd1292d OR matchd1291d;
	-- d1293d
	sted1293d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1293d,
			Enable=>Enabled1293d,
			match=>matchd1293d,
			run=>run);

	Enabled1293d <= matchd1292d;
	-- d1294d
	sted1294d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1294d,
			Enable=>Enabled1294d,
			match=>matchd1294d,
			run=>run);

	Enabled1294d <= matchd1293d OR matchd1294d;
	-- d1295d
	sted1295d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1295d,
			Enable=>Enabled1295d,
			match=>matchd1295d,
			run=>run);

	Enabled1295d <= matchd1294d;
	-- d1296d
	sted1296d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1296d,
			Enable=>Enabled1296d,
			match=>matchd1296d,
			run=>run);

	Enabled1296d <= matchd1295d;
	-- d1297d
	sted1297d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1297d,
			Enable=>Enabled1297d,
			match=>matchd1297d,
			run=>run);

	Enabled1297d <= matchd1296d;
	-- d1298d
	sted1298d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1298d,
			Enable=>Enabled1298d,
			match=>matchd1298d,
			run=>run);

	Enabled1298d <= matchd1297d;
	-- d1300d
	sted1300d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1300d,
			Enable=>Enabled1300d,
			match=>matchd1300d,
			run=>run);

	-- d1301d
	sted1301d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1301d,
			Enable=>Enabled1301d,
			match=>matchd1301d,
			run=>run);

	Enabled1301d <= matchd1300d;
	-- d1302d
	sted1302d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1302d,
			Enable=>Enabled1302d,
			match=>matchd1302d,
			run=>run);

	Enabled1302d <= matchd1301d;
	-- d1303d
	sted1303d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1303d,
			Enable=>Enabled1303d,
			match=>matchd1303d,
			run=>run);

	Enabled1303d <= matchd1302d;
	-- d1304d
	sted1304d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1304d,
			Enable=>Enabled1304d,
			match=>matchd1304d,
			run=>run);

	Enabled1304d <= matchd1303d;
	-- d1305d
	sted1305d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1305d,
			Enable=>Enabled1305d,
			match=>matchd1305d,
			run=>run);

	Enabled1305d <= matchd1305d OR matchd1304d;
	-- d1306d
	sted1306d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1306d,
			Enable=>Enabled1306d,
			match=>matchd1306d,
			run=>run);

	Enabled1306d <= matchd1305d;
	-- d1307d
	sted1307d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1307d,
			Enable=>Enabled1307d,
			match=>matchd1307d,
			run=>run);

	Enabled1307d <= matchd1306d OR matchd1307d;
	-- d1308d
	sted1308d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1308d,
			Enable=>Enabled1308d,
			match=>matchd1308d,
			run=>run);

	Enabled1308d <= matchd1307d;
	-- d1309d
	sted1309d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1309d,
			Enable=>Enabled1309d,
			match=>matchd1309d,
			run=>run);

	Enabled1309d <= matchd1308d;
	-- d1310d
	sted1310d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1310d,
			Enable=>Enabled1310d,
			match=>matchd1310d,
			run=>run);

	Enabled1310d <= matchd1309d;
	-- d1311d
	sted1311d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1311d,
			Enable=>Enabled1311d,
			match=>matchd1311d,
			run=>run);

	Enabled1311d <= matchd1310d;
	-- d1312d
	sted1312d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1312d,
			Enable=>Enabled1312d,
			match=>matchd1312d,
			run=>run);

	reports(58) <= matchd1312d;
	Enabled1312d <= matchd1311d;
	-- d1313d
	sted1313d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1313d,
			Enable=>Enabled1313d,
			match=>matchd1313d,
			run=>run);

	-- d1314d
	sted1314d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1314d,
			Enable=>Enabled1314d,
			match=>matchd1314d,
			run=>run);

	Enabled1314d <= matchd1314d OR matchd1313d;
	-- d1315d
	sted1315d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1315d,
			Enable=>Enabled1315d,
			match=>matchd1315d,
			run=>run);

	Enabled1315d <= matchd1314d;
	-- d1316d
	sted1316d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1316d,
			Enable=>Enabled1316d,
			match=>matchd1316d,
			run=>run);

	Enabled1316d <= matchd1315d;
	-- d1317d
	sted1317d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1317d,
			Enable=>Enabled1317d,
			match=>matchd1317d,
			run=>run);

	Enabled1317d <= matchd1316d;
	-- d1318d
	sted1318d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1318d,
			Enable=>Enabled1318d,
			match=>matchd1318d,
			run=>run);

	Enabled1318d <= matchd1317d;
	-- d1319d
	sted1319d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1319d,
			Enable=>Enabled1319d,
			match=>matchd1319d,
			run=>run);

	Enabled1319d <= matchd1318d;
	-- d1320d
	sted1320d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1320d,
			Enable=>Enabled1320d,
			match=>matchd1320d,
			run=>run);

	Enabled1320d <= matchd1320d OR matchd1319d;
	-- d1321d
	sted1321d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1321d,
			Enable=>Enabled1321d,
			match=>matchd1321d,
			run=>run);

	Enabled1321d <= matchd1320d;
	-- d1322d
	sted1322d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1322d,
			Enable=>Enabled1322d,
			match=>matchd1322d,
			run=>run);

	Enabled1322d <= matchd1321d;
	-- d1323d
	sted1323d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1323d,
			Enable=>Enabled1323d,
			match=>matchd1323d,
			run=>run);

	Enabled1323d <= matchd1322d;
	-- d1324d
	sted1324d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1324d,
			Enable=>Enabled1324d,
			match=>matchd1324d,
			run=>run);

	Enabled1324d <= matchd1323d;
	-- d1325d
	sted1325d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1325d,
			Enable=>Enabled1325d,
			match=>matchd1325d,
			run=>run);

	Enabled1325d <= matchd1324d OR matchd1325d;
	-- d1326d
	sted1326d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1326d,
			Enable=>Enabled1326d,
			match=>matchd1326d,
			run=>run);

	Enabled1326d <= matchd1325d;
	-- d1327d
	sted1327d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1327d,
			Enable=>Enabled1327d,
			match=>matchd1327d,
			run=>run);

	Enabled1327d <= matchd1326d;
	-- d1328d
	sted1328d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1328d,
			Enable=>Enabled1328d,
			match=>matchd1328d,
			run=>run);

	Enabled1328d <= matchd1327d;
	-- d1329d
	sted1329d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1329d,
			Enable=>Enabled1329d,
			match=>matchd1329d,
			run=>run);

	Enabled1329d <= matchd1328d;
	-- d1330d
	sted1330d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1330d,
			Enable=>Enabled1330d,
			match=>matchd1330d,
			run=>run);

	reports(59) <= matchd1330d;
	Enabled1330d <= matchd1329d;
	-- d1331d
	sted1331d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1331d,
			Enable=>Enabled1331d,
			match=>matchd1331d,
			run=>run);

	-- d1332d
	sted1332d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1332d,
			Enable=>Enabled1332d,
			match=>matchd1332d,
			run=>run);

	Enabled1332d <= matchd1332d OR matchd1331d;
	-- d1333d
	sted1333d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1333d,
			Enable=>Enabled1333d,
			match=>matchd1333d,
			run=>run);

	Enabled1333d <= matchd1332d;
	-- d1334d
	sted1334d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1334d,
			Enable=>Enabled1334d,
			match=>matchd1334d,
			run=>run);

	Enabled1334d <= matchd1333d;
	-- d1335d
	sted1335d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1335d,
			Enable=>Enabled1335d,
			match=>matchd1335d,
			run=>run);

	Enabled1335d <= matchd1334d;
	-- d1336d
	sted1336d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1336d,
			Enable=>Enabled1336d,
			match=>matchd1336d,
			run=>run);

	Enabled1336d <= matchd1335d;
	-- d1337d
	sted1337d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1337d,
			Enable=>Enabled1337d,
			match=>matchd1337d,
			run=>run);

	Enabled1337d <= matchd1337d OR matchd1336d;
	-- d1338d
	sted1338d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1338d,
			Enable=>Enabled1338d,
			match=>matchd1338d,
			run=>run);

	Enabled1338d <= matchd1337d;
	-- d1339d
	sted1339d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1339d,
			Enable=>Enabled1339d,
			match=>matchd1339d,
			run=>run);

	Enabled1339d <= matchd1338d;
	-- d1340d
	sted1340d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1340d,
			Enable=>Enabled1340d,
			match=>matchd1340d,
			run=>run);

	Enabled1340d <= matchd1339d;
	-- d1341d
	sted1341d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1341d,
			Enable=>Enabled1341d,
			match=>matchd1341d,
			run=>run);

	Enabled1341d <= matchd1340d;
	-- d1342d
	sted1342d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1342d,
			Enable=>Enabled1342d,
			match=>matchd1342d,
			run=>run);

	Enabled1342d <= matchd1341d OR matchd1342d;
	-- d1343d
	sted1343d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1343d,
			Enable=>Enabled1343d,
			match=>matchd1343d,
			run=>run);

	Enabled1343d <= matchd1342d;
	-- d1344d
	sted1344d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1344d,
			Enable=>Enabled1344d,
			match=>matchd1344d,
			run=>run);

	Enabled1344d <= matchd1343d;
	-- d1345d
	sted1345d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1345d,
			Enable=>Enabled1345d,
			match=>matchd1345d,
			run=>run);

	Enabled1345d <= matchd1344d;
	-- d1346d
	sted1346d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1346d,
			Enable=>Enabled1346d,
			match=>matchd1346d,
			run=>run);

	reports(60) <= matchd1346d;
	Enabled1346d <= matchd1345d;
	-- d1347d
	sted1347d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1347d,
			Enable=>Enabled1347d,
			match=>matchd1347d,
			run=>run);

	-- d1348d
	sted1348d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1348d,
			Enable=>Enabled1348d,
			match=>matchd1348d,
			run=>run);

	Enabled1348d <= matchd1348d OR matchd1347d;
	-- d1349d
	sted1349d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1349d,
			Enable=>Enabled1349d,
			match=>matchd1349d,
			run=>run);

	Enabled1349d <= matchd1348d;
	-- d1350d
	sted1350d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1350d,
			Enable=>Enabled1350d,
			match=>matchd1350d,
			run=>run);

	Enabled1350d <= matchd1349d;
	-- d1351d
	sted1351d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1351d,
			Enable=>Enabled1351d,
			match=>matchd1351d,
			run=>run);

	Enabled1351d <= matchd1350d;
	-- d1352d
	sted1352d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1352d,
			Enable=>Enabled1352d,
			match=>matchd1352d,
			run=>run);

	Enabled1352d <= matchd1351d;
	-- d1353d
	sted1353d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1353d,
			Enable=>Enabled1353d,
			match=>matchd1353d,
			run=>run);

	Enabled1353d <= matchd1353d OR matchd1352d;
	-- d1354d
	sted1354d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1354d,
			Enable=>Enabled1354d,
			match=>matchd1354d,
			run=>run);

	Enabled1354d <= matchd1353d;
	-- d1355d
	sted1355d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1355d,
			Enable=>Enabled1355d,
			match=>matchd1355d,
			run=>run);

	Enabled1355d <= matchd1354d;
	-- d1356d
	sted1356d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1356d,
			Enable=>Enabled1356d,
			match=>matchd1356d,
			run=>run);

	Enabled1356d <= matchd1355d;
	-- d1357d
	sted1357d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1357d,
			Enable=>Enabled1357d,
			match=>matchd1357d,
			run=>run);

	Enabled1357d <= matchd1356d;
	-- d1358d
	sted1358d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1358d,
			Enable=>Enabled1358d,
			match=>matchd1358d,
			run=>run);

	reports(61) <= matchd1358d;
	Enabled1358d <= matchd1357d;
	-- d1359d
	sted1359d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1359d,
			Enable=>Enabled1359d,
			match=>matchd1359d,
			run=>run);

	-- d1360d
	sted1360d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1360d,
			Enable=>Enabled1360d,
			match=>matchd1360d,
			run=>run);

	Enabled1360d <= matchd1359d OR matchd1360d;
	-- d1361d
	sted1361d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1361d,
			Enable=>Enabled1361d,
			match=>matchd1361d,
			run=>run);

	Enabled1361d <= matchd1360d;
	-- d1362d
	sted1362d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1362d,
			Enable=>Enabled1362d,
			match=>matchd1362d,
			run=>run);

	Enabled1362d <= matchd1361d;
	-- d1363d
	sted1363d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1363d,
			Enable=>Enabled1363d,
			match=>matchd1363d,
			run=>run);

	Enabled1363d <= matchd1362d;
	-- d1364d
	sted1364d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1364d,
			Enable=>Enabled1364d,
			match=>matchd1364d,
			run=>run);

	Enabled1364d <= matchd1363d;
	-- d1365d
	sted1365d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1365d,
			Enable=>Enabled1365d,
			match=>matchd1365d,
			run=>run);

	Enabled1365d <= matchd1364d;
	-- d1366d
	sted1366d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1366d,
			Enable=>Enabled1366d,
			match=>matchd1366d,
			run=>run);

	Enabled1366d <= matchd1366d OR matchd1365d;
	-- d1367d
	sted1367d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1367d,
			Enable=>Enabled1367d,
			match=>matchd1367d,
			run=>run);

	Enabled1367d <= matchd1366d;
	-- d1368d
	sted1368d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1368d,
			Enable=>Enabled1368d,
			match=>matchd1368d,
			run=>run);

	Enabled1368d <= matchd1367d;
	-- d1369d
	sted1369d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1369d,
			Enable=>Enabled1369d,
			match=>matchd1369d,
			run=>run);

	Enabled1369d <= matchd1368d;
	-- d1370d
	sted1370d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1370d,
			Enable=>Enabled1370d,
			match=>matchd1370d,
			run=>run);

	Enabled1370d <= matchd1369d;
	-- d1371d
	sted1371d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1371d,
			Enable=>Enabled1371d,
			match=>matchd1371d,
			run=>run);

	Enabled1371d <= matchd1371d OR matchd1370d;
	-- d1372d
	sted1372d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1372d,
			Enable=>Enabled1372d,
			match=>matchd1372d,
			run=>run);

	Enabled1372d <= matchd1371d;
	-- d1373d
	sted1373d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1373d,
			Enable=>Enabled1373d,
			match=>matchd1373d,
			run=>run);

	Enabled1373d <= matchd1372d;
	-- d1374d
	sted1374d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1374d,
			Enable=>Enabled1374d,
			match=>matchd1374d,
			run=>run);

	Enabled1374d <= matchd1373d;
	-- d1375d
	sted1375d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1375d,
			Enable=>Enabled1375d,
			match=>matchd1375d,
			run=>run);

	Enabled1375d <= matchd1374d;
	-- d1376d
	sted1376d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1376d,
			Enable=>Enabled1376d,
			match=>matchd1376d,
			run=>run);

	reports(62) <= matchd1376d;
	Enabled1376d <= matchd1375d;
	-- d1377d
	sted1377d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1377d,
			Enable=>Enabled1377d,
			match=>matchd1377d,
			run=>run);

	-- d1378d
	sted1378d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1378d,
			Enable=>Enabled1378d,
			match=>matchd1378d,
			run=>run);

	Enabled1378d <= matchd1377d OR matchd1378d;
	-- d1379d
	sted1379d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1379d,
			Enable=>Enabled1379d,
			match=>matchd1379d,
			run=>run);

	Enabled1379d <= matchd1378d;
	-- d1380d
	sted1380d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1380d,
			Enable=>Enabled1380d,
			match=>matchd1380d,
			run=>run);

	Enabled1380d <= matchd1379d;
	-- d1381d
	sted1381d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1381d,
			Enable=>Enabled1381d,
			match=>matchd1381d,
			run=>run);

	Enabled1381d <= matchd1380d;
	-- d1382d
	sted1382d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1382d,
			Enable=>Enabled1382d,
			match=>matchd1382d,
			run=>run);

	Enabled1382d <= matchd1381d;
	-- d1383d
	sted1383d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1383d,
			Enable=>Enabled1383d,
			match=>matchd1383d,
			run=>run);

	Enabled1383d <= matchd1382d OR matchd1383d;
	-- d1384d
	sted1384d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1384d,
			Enable=>Enabled1384d,
			match=>matchd1384d,
			run=>run);

	Enabled1384d <= matchd1383d;
	-- d1385d
	sted1385d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1385d,
			Enable=>Enabled1385d,
			match=>matchd1385d,
			run=>run);

	Enabled1385d <= matchd1384d;
	-- d1386d
	sted1386d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1386d,
			Enable=>Enabled1386d,
			match=>matchd1386d,
			run=>run);

	reports(63) <= matchd1386d;
	Enabled1386d <= matchd1385d;
	-- d1387d
	sted1387d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1387d,
			Enable=>Enabled1387d,
			match=>matchd1387d,
			run=>run);

	-- d1388d
	sted1388d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1388d,
			Enable=>Enabled1388d,
			match=>matchd1388d,
			run=>run);

	Enabled1388d <= matchd1387d OR matchd1388d;
	-- d1389d
	sted1389d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1389d,
			Enable=>Enabled1389d,
			match=>matchd1389d,
			run=>run);

	Enabled1389d <= matchd1388d;
	-- d1390d
	sted1390d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1390d,
			Enable=>Enabled1390d,
			match=>matchd1390d,
			run=>run);

	Enabled1390d <= matchd1389d;
	-- d1391d
	sted1391d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1391d,
			Enable=>Enabled1391d,
			match=>matchd1391d,
			run=>run);

	Enabled1391d <= matchd1390d;
	-- d1392d
	sted1392d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1392d,
			Enable=>Enabled1392d,
			match=>matchd1392d,
			run=>run);

	Enabled1392d <= matchd1392d OR matchd1391d;
	-- d1393d
	sted1393d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1393d,
			Enable=>Enabled1393d,
			match=>matchd1393d,
			run=>run);

	Enabled1393d <= matchd1392d;
	-- d1394d
	sted1394d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1394d,
			Enable=>Enabled1394d,
			match=>matchd1394d,
			run=>run);

	Enabled1394d <= matchd1393d;
	-- d1395d
	sted1395d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1395d,
			Enable=>Enabled1395d,
			match=>matchd1395d,
			run=>run);

	Enabled1395d <= matchd1394d;
	-- d1396d
	sted1396d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1396d,
			Enable=>Enabled1396d,
			match=>matchd1396d,
			run=>run);

	Enabled1396d <= matchd1395d;
	-- d1397d
	sted1397d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1397d,
			Enable=>Enabled1397d,
			match=>matchd1397d,
			run=>run);

	Enabled1397d <= matchd1396d;
	-- d1398d
	sted1398d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1398d,
			Enable=>Enabled1398d,
			match=>matchd1398d,
			run=>run);

	Enabled1398d <= matchd1397d OR matchd1398d;
	-- d1399d
	sted1399d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1399d,
			Enable=>Enabled1399d,
			match=>matchd1399d,
			run=>run);

	Enabled1399d <= matchd1398d;
	-- d1400d
	sted1400d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1400d,
			Enable=>Enabled1400d,
			match=>matchd1400d,
			run=>run);

	Enabled1400d <= matchd1399d;
	-- d1401d
	sted1401d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1401d,
			Enable=>Enabled1401d,
			match=>matchd1401d,
			run=>run);

	Enabled1401d <= matchd1400d;
	-- d1402d
	sted1402d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1402d,
			Enable=>Enabled1402d,
			match=>matchd1402d,
			run=>run);

	reports(64) <= matchd1402d;
	Enabled1402d <= matchd1401d;
	-- d1403d
	sted1403d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1403d,
			Enable=>Enabled1403d,
			match=>matchd1403d,
			run=>run);

	-- d1404d
	sted1404d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1404d,
			Enable=>Enabled1404d,
			match=>matchd1404d,
			run=>run);

	Enabled1404d <= matchd1404d OR matchd1403d;
	-- d1405d
	sted1405d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1405d,
			Enable=>Enabled1405d,
			match=>matchd1405d,
			run=>run);

	Enabled1405d <= matchd1404d;
	-- d1406d
	sted1406d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1406d,
			Enable=>Enabled1406d,
			match=>matchd1406d,
			run=>run);

	Enabled1406d <= matchd1405d;
	-- d1407d
	sted1407d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1407d,
			Enable=>Enabled1407d,
			match=>matchd1407d,
			run=>run);

	Enabled1407d <= matchd1406d;
	-- d1408d
	sted1408d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1408d,
			Enable=>Enabled1408d,
			match=>matchd1408d,
			run=>run);

	Enabled1408d <= matchd1407d;
	-- d1409d
	sted1409d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1409d,
			Enable=>Enabled1409d,
			match=>matchd1409d,
			run=>run);

	Enabled1409d <= matchd1409d OR matchd1408d;
	-- d1410d
	sted1410d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1410d,
			Enable=>Enabled1410d,
			match=>matchd1410d,
			run=>run);

	Enabled1410d <= matchd1409d;
	-- d1411d
	sted1411d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1411d,
			Enable=>Enabled1411d,
			match=>matchd1411d,
			run=>run);

	Enabled1411d <= matchd1410d;
	-- d1412d
	sted1412d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1412d,
			Enable=>Enabled1412d,
			match=>matchd1412d,
			run=>run);

	Enabled1412d <= matchd1411d;
	-- d1413d
	sted1413d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1413d,
			Enable=>Enabled1413d,
			match=>matchd1413d,
			run=>run);

	reports(65) <= matchd1413d;
	Enabled1413d <= matchd1412d;
	-- d1414d
	sted1414d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1414d,
			Enable=>Enabled1414d,
			match=>matchd1414d,
			run=>run);

	-- d1415d
	sted1415d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1415d,
			Enable=>Enabled1415d,
			match=>matchd1415d,
			run=>run);

	Enabled1415d <= matchd1414d OR matchd1415d;
	-- d1416d
	sted1416d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1416d,
			Enable=>Enabled1416d,
			match=>matchd1416d,
			run=>run);

	Enabled1416d <= matchd1415d;
	-- d1417d
	sted1417d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1417d,
			Enable=>Enabled1417d,
			match=>matchd1417d,
			run=>run);

	Enabled1417d <= matchd1416d;
	-- d1418d
	sted1418d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1418d,
			Enable=>Enabled1418d,
			match=>matchd1418d,
			run=>run);

	Enabled1418d <= matchd1417d;
	-- d1419d
	sted1419d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1419d,
			Enable=>Enabled1419d,
			match=>matchd1419d,
			run=>run);

	Enabled1419d <= matchd1418d;
	-- d1420d
	sted1420d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1420d,
			Enable=>Enabled1420d,
			match=>matchd1420d,
			run=>run);

	Enabled1420d <= matchd1420d OR matchd1419d;
	-- d1421d
	sted1421d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1421d,
			Enable=>Enabled1421d,
			match=>matchd1421d,
			run=>run);

	Enabled1421d <= matchd1420d;
	-- d1422d
	sted1422d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1422d,
			Enable=>Enabled1422d,
			match=>matchd1422d,
			run=>run);

	Enabled1422d <= matchd1421d;
	-- d1423d
	sted1423d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1423d,
			Enable=>Enabled1423d,
			match=>matchd1423d,
			run=>run);

	Enabled1423d <= matchd1422d;
	-- d1424d
	sted1424d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1424d,
			Enable=>Enabled1424d,
			match=>matchd1424d,
			run=>run);

	Enabled1424d <= matchd1423d;
	-- d1425d
	sted1425d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1425d,
			Enable=>Enabled1425d,
			match=>matchd1425d,
			run=>run);

	Enabled1425d <= matchd1425d OR matchd1424d;
	-- d1426d
	sted1426d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1426d,
			Enable=>Enabled1426d,
			match=>matchd1426d,
			run=>run);

	Enabled1426d <= matchd1425d;
	-- d1427d
	sted1427d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1427d,
			Enable=>Enabled1427d,
			match=>matchd1427d,
			run=>run);

	Enabled1427d <= matchd1426d;
	-- d1428d
	sted1428d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1428d,
			Enable=>Enabled1428d,
			match=>matchd1428d,
			run=>run);

	Enabled1428d <= matchd1427d;
	-- d1429d
	sted1429d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1429d,
			Enable=>Enabled1429d,
			match=>matchd1429d,
			run=>run);

	reports(66) <= matchd1429d;
	Enabled1429d <= matchd1428d;
	-- d1430d
	sted1430d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1430d,
			Enable=>Enabled1430d,
			match=>matchd1430d,
			run=>run);

	-- d1431d
	sted1431d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1431d,
			Enable=>Enabled1431d,
			match=>matchd1431d,
			run=>run);

	Enabled1431d <= matchd1431d OR matchd1430d;
	-- d1432d
	sted1432d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1432d,
			Enable=>Enabled1432d,
			match=>matchd1432d,
			run=>run);

	Enabled1432d <= matchd1431d;
	-- d1433d
	sted1433d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1433d,
			Enable=>Enabled1433d,
			match=>matchd1433d,
			run=>run);

	Enabled1433d <= matchd1432d;
	-- d1434d
	sted1434d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1434d,
			Enable=>Enabled1434d,
			match=>matchd1434d,
			run=>run);

	Enabled1434d <= matchd1433d;
	-- d1435d
	sted1435d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1435d,
			Enable=>Enabled1435d,
			match=>matchd1435d,
			run=>run);

	Enabled1435d <= matchd1434d;
	-- d1436d
	sted1436d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1436d,
			Enable=>Enabled1436d,
			match=>matchd1436d,
			run=>run);

	Enabled1436d <= matchd1435d;
	-- d1437d
	sted1437d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1437d,
			Enable=>Enabled1437d,
			match=>matchd1437d,
			run=>run);

	Enabled1437d <= matchd1436d OR matchd1437d;
	-- d1438d
	sted1438d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1438d,
			Enable=>Enabled1438d,
			match=>matchd1438d,
			run=>run);

	Enabled1438d <= matchd1437d;
	-- d1439d
	sted1439d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1439d,
			Enable=>Enabled1439d,
			match=>matchd1439d,
			run=>run);

	Enabled1439d <= matchd1438d;
	-- d1440d
	sted1440d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1440d,
			Enable=>Enabled1440d,
			match=>matchd1440d,
			run=>run);

	Enabled1440d <= matchd1439d;
	-- d1441d
	sted1441d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1441d,
			Enable=>Enabled1441d,
			match=>matchd1441d,
			run=>run);

	Enabled1441d <= matchd1440d;
	-- d1442d
	sted1442d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1442d,
			Enable=>Enabled1442d,
			match=>matchd1442d,
			run=>run);

	reports(67) <= matchd1442d;
	Enabled1442d <= matchd1441d;
	-- d1443d
	sted1443d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1443d,
			Enable=>Enabled1443d,
			match=>matchd1443d,
			run=>run);

	-- d1444d
	sted1444d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1444d,
			Enable=>Enabled1444d,
			match=>matchd1444d,
			run=>run);

	Enabled1444d <= matchd1444d OR matchd1443d;
	-- d1445d
	sted1445d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1445d,
			Enable=>Enabled1445d,
			match=>matchd1445d,
			run=>run);

	Enabled1445d <= matchd1444d;
	-- d1446d
	sted1446d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1446d,
			Enable=>Enabled1446d,
			match=>matchd1446d,
			run=>run);

	Enabled1446d <= matchd1445d;
	-- d1447d
	sted1447d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1447d,
			Enable=>Enabled1447d,
			match=>matchd1447d,
			run=>run);

	Enabled1447d <= matchd1446d;
	-- d1448d
	sted1448d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1448d,
			Enable=>Enabled1448d,
			match=>matchd1448d,
			run=>run);

	Enabled1448d <= matchd1447d;
	-- d1449d
	sted1449d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1449d,
			Enable=>Enabled1449d,
			match=>matchd1449d,
			run=>run);

	Enabled1449d <= matchd1449d OR matchd1448d;
	-- d1450d
	sted1450d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1450d,
			Enable=>Enabled1450d,
			match=>matchd1450d,
			run=>run);

	Enabled1450d <= matchd1449d;
	-- d1451d
	sted1451d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1451d,
			Enable=>Enabled1451d,
			match=>matchd1451d,
			run=>run);

	Enabled1451d <= matchd1450d;
	-- d1452d
	sted1452d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1452d,
			Enable=>Enabled1452d,
			match=>matchd1452d,
			run=>run);

	Enabled1452d <= matchd1451d;
	-- d1453d
	sted1453d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1453d,
			Enable=>Enabled1453d,
			match=>matchd1453d,
			run=>run);

	Enabled1453d <= matchd1452d;
	-- d1454d
	sted1454d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1454d,
			Enable=>Enabled1454d,
			match=>matchd1454d,
			run=>run);

	reports(68) <= matchd1454d;
	Enabled1454d <= matchd1453d;
	-- d1455d
	sted1455d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1455d,
			Enable=>Enabled1455d,
			match=>matchd1455d,
			run=>run);

	-- d1456d
	sted1456d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1456d,
			Enable=>Enabled1456d,
			match=>matchd1456d,
			run=>run);

	Enabled1456d <= matchd1455d OR matchd1456d;
	-- d1457d
	sted1457d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1457d,
			Enable=>Enabled1457d,
			match=>matchd1457d,
			run=>run);

	Enabled1457d <= matchd1456d;
	-- d1458d
	sted1458d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1458d,
			Enable=>Enabled1458d,
			match=>matchd1458d,
			run=>run);

	Enabled1458d <= matchd1457d;
	-- d1459d
	sted1459d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1459d,
			Enable=>Enabled1459d,
			match=>matchd1459d,
			run=>run);

	Enabled1459d <= matchd1458d;
	-- d1460d
	sted1460d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1460d,
			Enable=>Enabled1460d,
			match=>matchd1460d,
			run=>run);

	Enabled1460d <= matchd1459d;
	-- d1461d
	sted1461d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1461d,
			Enable=>Enabled1461d,
			match=>matchd1461d,
			run=>run);

	Enabled1461d <= matchd1460d;
	-- d1462d
	sted1462d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1462d,
			Enable=>Enabled1462d,
			match=>matchd1462d,
			run=>run);

	Enabled1462d <= matchd1461d;
	-- d1463d
	sted1463d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1463d,
			Enable=>Enabled1463d,
			match=>matchd1463d,
			run=>run);

	Enabled1463d <= matchd1463d OR matchd1462d;
	-- d1464d
	sted1464d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1464d,
			Enable=>Enabled1464d,
			match=>matchd1464d,
			run=>run);

	Enabled1464d <= matchd1463d;
	-- d1465d
	sted1465d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1465d,
			Enable=>Enabled1465d,
			match=>matchd1465d,
			run=>run);

	Enabled1465d <= matchd1464d;
	-- d1466d
	sted1466d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1466d,
			Enable=>Enabled1466d,
			match=>matchd1466d,
			run=>run);

	Enabled1466d <= matchd1465d;
	-- d1467d
	sted1467d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1467d,
			Enable=>Enabled1467d,
			match=>matchd1467d,
			run=>run);

	reports(69) <= matchd1467d;
	Enabled1467d <= matchd1466d;
	-- d1468d
	sted1468d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1468d,
			Enable=>Enabled1468d,
			match=>matchd1468d,
			run=>run);

	-- d1469d
	sted1469d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1469d,
			Enable=>Enabled1469d,
			match=>matchd1469d,
			run=>run);

	Enabled1469d <= matchd1469d OR matchd1468d;
	-- d1470d
	sted1470d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1470d,
			Enable=>Enabled1470d,
			match=>matchd1470d,
			run=>run);

	Enabled1470d <= matchd1469d;
	-- d1471d
	sted1471d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1471d,
			Enable=>Enabled1471d,
			match=>matchd1471d,
			run=>run);

	Enabled1471d <= matchd1470d;
	-- d1472d
	sted1472d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1472d,
			Enable=>Enabled1472d,
			match=>matchd1472d,
			run=>run);

	Enabled1472d <= matchd1471d;
	-- d1473d
	sted1473d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1473d,
			Enable=>Enabled1473d,
			match=>matchd1473d,
			run=>run);

	Enabled1473d <= matchd1472d;
	-- d1474d
	sted1474d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1474d,
			Enable=>Enabled1474d,
			match=>matchd1474d,
			run=>run);

	Enabled1474d <= matchd1473d;
	-- d1475d
	sted1475d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1475d,
			Enable=>Enabled1475d,
			match=>matchd1475d,
			run=>run);

	Enabled1475d <= matchd1474d OR matchd1475d;
	-- d1476d
	sted1476d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1476d,
			Enable=>Enabled1476d,
			match=>matchd1476d,
			run=>run);

	Enabled1476d <= matchd1475d;
	-- d1477d
	sted1477d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1477d,
			Enable=>Enabled1477d,
			match=>matchd1477d,
			run=>run);

	Enabled1477d <= matchd1476d;
	-- d1478d
	sted1478d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1478d,
			Enable=>Enabled1478d,
			match=>matchd1478d,
			run=>run);

	Enabled1478d <= matchd1477d;
	-- d1479d
	sted1479d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1479d,
			Enable=>Enabled1479d,
			match=>matchd1479d,
			run=>run);

	reports(70) <= matchd1479d;
	Enabled1479d <= matchd1478d;
	-- d1480d
	sted1480d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1480d,
			Enable=>Enabled1480d,
			match=>matchd1480d,
			run=>run);

	-- d1481d
	sted1481d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1481d,
			Enable=>Enabled1481d,
			match=>matchd1481d,
			run=>run);

	Enabled1481d <= matchd1481d OR matchd1480d;
	-- d1482d
	sted1482d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1482d,
			Enable=>Enabled1482d,
			match=>matchd1482d,
			run=>run);

	Enabled1482d <= matchd1481d;
	-- d1483d
	sted1483d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1483d,
			Enable=>Enabled1483d,
			match=>matchd1483d,
			run=>run);

	Enabled1483d <= matchd1482d;
	-- d1484d
	sted1484d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1484d,
			Enable=>Enabled1484d,
			match=>matchd1484d,
			run=>run);

	Enabled1484d <= matchd1483d;
	-- d1485d
	sted1485d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1485d,
			Enable=>Enabled1485d,
			match=>matchd1485d,
			run=>run);

	Enabled1485d <= matchd1484d;
	-- d1486d
	sted1486d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1486d,
			Enable=>Enabled1486d,
			match=>matchd1486d,
			run=>run);

	Enabled1486d <= matchd1485d;
	-- d1487d
	sted1487d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1487d,
			Enable=>Enabled1487d,
			match=>matchd1487d,
			run=>run);

	Enabled1487d <= matchd1486d;
	-- d1488d
	sted1488d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1488d,
			Enable=>Enabled1488d,
			match=>matchd1488d,
			run=>run);

	Enabled1488d <= matchd1487d OR matchd1488d;
	-- d1489d
	sted1489d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1489d,
			Enable=>Enabled1489d,
			match=>matchd1489d,
			run=>run);

	Enabled1489d <= matchd1488d;
	-- d1490d
	sted1490d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1490d,
			Enable=>Enabled1490d,
			match=>matchd1490d,
			run=>run);

	Enabled1490d <= matchd1489d;
	-- d1491d
	sted1491d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1491d,
			Enable=>Enabled1491d,
			match=>matchd1491d,
			run=>run);

	Enabled1491d <= matchd1490d;
	-- d1492d
	sted1492d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1492d,
			Enable=>Enabled1492d,
			match=>matchd1492d,
			run=>run);

	reports(71) <= matchd1492d;
	Enabled1492d <= matchd1491d;
	-- d1493d
	sted1493d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1493d,
			Enable=>Enabled1493d,
			match=>matchd1493d,
			run=>run);

	-- d1494d
	sted1494d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1494d,
			Enable=>Enabled1494d,
			match=>matchd1494d,
			run=>run);

	Enabled1494d <= matchd1493d OR matchd1494d;
	-- d1495d
	sted1495d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1495d,
			Enable=>Enabled1495d,
			match=>matchd1495d,
			run=>run);

	Enabled1495d <= matchd1494d;
	-- d1496d
	sted1496d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1496d,
			Enable=>Enabled1496d,
			match=>matchd1496d,
			run=>run);

	Enabled1496d <= matchd1495d;
	-- d1497d
	sted1497d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1497d,
			Enable=>Enabled1497d,
			match=>matchd1497d,
			run=>run);

	Enabled1497d <= matchd1496d;
	-- d1498d
	sted1498d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1498d,
			Enable=>Enabled1498d,
			match=>matchd1498d,
			run=>run);

	Enabled1498d <= matchd1497d;
	-- d1499d
	sted1499d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1499d,
			Enable=>Enabled1499d,
			match=>matchd1499d,
			run=>run);

	Enabled1499d <= matchd1498d;
	-- d1500d
	sted1500d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1500d,
			Enable=>Enabled1500d,
			match=>matchd1500d,
			run=>run);

	Enabled1500d <= matchd1500d OR matchd1499d;
	-- d1501d
	sted1501d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1501d,
			Enable=>Enabled1501d,
			match=>matchd1501d,
			run=>run);

	Enabled1501d <= matchd1500d;
	-- d1502d
	sted1502d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1502d,
			Enable=>Enabled1502d,
			match=>matchd1502d,
			run=>run);

	Enabled1502d <= matchd1501d;
	-- d1503d
	sted1503d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1503d,
			Enable=>Enabled1503d,
			match=>matchd1503d,
			run=>run);

	Enabled1503d <= matchd1502d;
	-- d1504d
	sted1504d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1504d,
			Enable=>Enabled1504d,
			match=>matchd1504d,
			run=>run);

	Enabled1504d <= matchd1503d;
	-- d1505d
	sted1505d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1505d,
			Enable=>Enabled1505d,
			match=>matchd1505d,
			run=>run);

	Enabled1505d <= matchd1504d OR matchd1505d;
	-- d1506d
	sted1506d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1506d,
			Enable=>Enabled1506d,
			match=>matchd1506d,
			run=>run);

	Enabled1506d <= matchd1505d;
	-- d1507d
	sted1507d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1507d,
			Enable=>Enabled1507d,
			match=>matchd1507d,
			run=>run);

	Enabled1507d <= matchd1506d;
	-- d1508d
	sted1508d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1508d,
			Enable=>Enabled1508d,
			match=>matchd1508d,
			run=>run);

	Enabled1508d <= matchd1507d;
	-- d1509d
	sted1509d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1509d,
			Enable=>Enabled1509d,
			match=>matchd1509d,
			run=>run);

	reports(72) <= matchd1509d;
	Enabled1509d <= matchd1508d;
	-- d1510d
	sted1510d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1510d,
			Enable=>Enabled1510d,
			match=>matchd1510d,
			run=>run);

	-- d1511d
	sted1511d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1511d,
			Enable=>Enabled1511d,
			match=>matchd1511d,
			run=>run);

	Enabled1511d <= matchd1511d OR matchd1510d;
	-- d1512d
	sted1512d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1512d,
			Enable=>Enabled1512d,
			match=>matchd1512d,
			run=>run);

	Enabled1512d <= matchd1511d;
	-- d1513d
	sted1513d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1513d,
			Enable=>Enabled1513d,
			match=>matchd1513d,
			run=>run);

	Enabled1513d <= matchd1512d;
	-- d1514d
	sted1514d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1514d,
			Enable=>Enabled1514d,
			match=>matchd1514d,
			run=>run);

	Enabled1514d <= matchd1513d;
	-- d1515d
	sted1515d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1515d,
			Enable=>Enabled1515d,
			match=>matchd1515d,
			run=>run);

	Enabled1515d <= matchd1514d;
	-- d1516d
	sted1516d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1516d,
			Enable=>Enabled1516d,
			match=>matchd1516d,
			run=>run);

	Enabled1516d <= matchd1516d OR matchd1515d;
	-- d1517d
	sted1517d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1517d,
			Enable=>Enabled1517d,
			match=>matchd1517d,
			run=>run);

	Enabled1517d <= matchd1516d;
	-- d1518d
	sted1518d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1518d,
			Enable=>Enabled1518d,
			match=>matchd1518d,
			run=>run);

	Enabled1518d <= matchd1517d;
	-- d1519d
	sted1519d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1519d,
			Enable=>Enabled1519d,
			match=>matchd1519d,
			run=>run);

	Enabled1519d <= matchd1518d;
	-- d1520d
	sted1520d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1520d,
			Enable=>Enabled1520d,
			match=>matchd1520d,
			run=>run);

	Enabled1520d <= matchd1519d;
	-- d1521d
	sted1521d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1521d,
			Enable=>Enabled1521d,
			match=>matchd1521d,
			run=>run);

	Enabled1521d <= matchd1520d;
	-- d1522d
	sted1522d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1522d,
			Enable=>Enabled1522d,
			match=>matchd1522d,
			run=>run);

	Enabled1522d <= matchd1521d OR matchd1522d;
	-- d1523d
	sted1523d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1523d,
			Enable=>Enabled1523d,
			match=>matchd1523d,
			run=>run);

	Enabled1523d <= matchd1522d;
	-- d1524d
	sted1524d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1524d,
			Enable=>Enabled1524d,
			match=>matchd1524d,
			run=>run);

	Enabled1524d <= matchd1523d;
	-- d1525d
	sted1525d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1525d,
			Enable=>Enabled1525d,
			match=>matchd1525d,
			run=>run);

	Enabled1525d <= matchd1524d;
	-- d1526d
	sted1526d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1526d,
			Enable=>Enabled1526d,
			match=>matchd1526d,
			run=>run);

	reports(73) <= matchd1526d;
	Enabled1526d <= matchd1525d;
	-- d1527d
	sted1527d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1527d,
			Enable=>Enabled1527d,
			match=>matchd1527d,
			run=>run);

	-- d1528d
	sted1528d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1528d,
			Enable=>Enabled1528d,
			match=>matchd1528d,
			run=>run);

	Enabled1528d <= matchd1527d;
	-- d1529d
	sted1529d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1529d,
			Enable=>Enabled1529d,
			match=>matchd1529d,
			run=>run);

	Enabled1529d <= matchd1528d;
	-- d1530d
	sted1530d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1530d,
			Enable=>Enabled1530d,
			match=>matchd1530d,
			run=>run);

	Enabled1530d <= matchd1529d;
	-- d1531d
	sted1531d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1531d,
			Enable=>Enabled1531d,
			match=>matchd1531d,
			run=>run);

	Enabled1531d <= matchd1530d;
	-- d1532d
	sted1532d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1532d,
			Enable=>Enabled1532d,
			match=>matchd1532d,
			run=>run);

	Enabled1532d <= matchd1531d;
	-- d1533d
	sted1533d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1533d,
			Enable=>Enabled1533d,
			match=>matchd1533d,
			run=>run);

	Enabled1533d <= matchd1532d;
	-- d1534d
	sted1534d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1534d,
			Enable=>Enabled1534d,
			match=>matchd1534d,
			run=>run);

	Enabled1534d <= matchd1533d;
	-- d1535d
	sted1535d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1535d,
			Enable=>Enabled1535d,
			match=>matchd1535d,
			run=>run);

	Enabled1535d <= matchd1534d;
	-- d1536d
	sted1536d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1536d,
			Enable=>Enabled1536d,
			match=>matchd1536d,
			run=>run);

	Enabled1536d <= matchd1535d;
	-- d1537d
	sted1537d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1537d,
			Enable=>Enabled1537d,
			match=>matchd1537d,
			run=>run);

	Enabled1537d <= matchd1537d OR matchd1536d;
	-- d1538d
	sted1538d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1538d,
			Enable=>Enabled1538d,
			match=>matchd1538d,
			run=>run);

	Enabled1538d <= matchd1537d;
	-- d1539d
	sted1539d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1539d,
			Enable=>Enabled1539d,
			match=>matchd1539d,
			run=>run);

	Enabled1539d <= matchd1538d;
	-- d1540d
	sted1540d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1540d,
			Enable=>Enabled1540d,
			match=>matchd1540d,
			run=>run);

	Enabled1540d <= matchd1539d;
	-- d1541d
	sted1541d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1541d,
			Enable=>Enabled1541d,
			match=>matchd1541d,
			run=>run);

	reports(74) <= matchd1541d;
	Enabled1541d <= matchd1540d;
	-- d1542d
	sted1542d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1542d,
			Enable=>Enabled1542d,
			match=>matchd1542d,
			run=>run);

	-- d1543d
	sted1543d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1543d,
			Enable=>Enabled1543d,
			match=>matchd1543d,
			run=>run);

	Enabled1543d <= matchd1542d;
	-- d1544d
	sted1544d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1544d,
			Enable=>Enabled1544d,
			match=>matchd1544d,
			run=>run);

	Enabled1544d <= matchd1543d;
	-- d1545d
	sted1545d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1545d,
			Enable=>Enabled1545d,
			match=>matchd1545d,
			run=>run);

	Enabled1545d <= matchd1544d;
	-- d1546d
	sted1546d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1546d,
			Enable=>Enabled1546d,
			match=>matchd1546d,
			run=>run);

	Enabled1546d <= matchd1545d;
	-- d1547d
	sted1547d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1547d,
			Enable=>Enabled1547d,
			match=>matchd1547d,
			run=>run);

	Enabled1547d <= matchd1546d;
	-- d1548d
	sted1548d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1548d,
			Enable=>Enabled1548d,
			match=>matchd1548d,
			run=>run);

	Enabled1548d <= matchd1548d OR matchd1547d;
	-- d1549d
	sted1549d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1549d,
			Enable=>Enabled1549d,
			match=>matchd1549d,
			run=>run);

	Enabled1549d <= matchd1548d;
	-- d1550d
	sted1550d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1550d,
			Enable=>Enabled1550d,
			match=>matchd1550d,
			run=>run);

	Enabled1550d <= matchd1550d OR matchd1549d;
	-- d1551d
	sted1551d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1551d,
			Enable=>Enabled1551d,
			match=>matchd1551d,
			run=>run);

	Enabled1551d <= matchd1550d;
	-- d1552d
	sted1552d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1552d,
			Enable=>Enabled1552d,
			match=>matchd1552d,
			run=>run);

	Enabled1552d <= matchd1551d;
	-- d1553d
	sted1553d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1553d,
			Enable=>Enabled1553d,
			match=>matchd1553d,
			run=>run);

	Enabled1553d <= matchd1552d;
	-- d1554d
	sted1554d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1554d,
			Enable=>Enabled1554d,
			match=>matchd1554d,
			run=>run);

	Enabled1554d <= matchd1553d;
	-- d1555d
	sted1555d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1555d,
			Enable=>Enabled1555d,
			match=>matchd1555d,
			run=>run);

	reports(75) <= matchd1555d;
	Enabled1555d <= matchd1554d;
	-- d1556d
	sted1556d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1556d,
			Enable=>Enabled1556d,
			match=>matchd1556d,
			run=>run);

	-- d1557d
	sted1557d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1557d,
			Enable=>Enabled1557d,
			match=>matchd1557d,
			run=>run);

	Enabled1557d <= matchd1557d OR matchd1556d;
	-- d1558d
	sted1558d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1558d,
			Enable=>Enabled1558d,
			match=>matchd1558d,
			run=>run);

	Enabled1558d <= matchd1557d;
	-- d1559d
	sted1559d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1559d,
			Enable=>Enabled1559d,
			match=>matchd1559d,
			run=>run);

	Enabled1559d <= matchd1558d;
	-- d1560d
	sted1560d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1560d,
			Enable=>Enabled1560d,
			match=>matchd1560d,
			run=>run);

	Enabled1560d <= matchd1559d;
	-- d1561d
	sted1561d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1561d,
			Enable=>Enabled1561d,
			match=>matchd1561d,
			run=>run);

	Enabled1561d <= matchd1560d;
	-- d1562d
	sted1562d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1562d,
			Enable=>Enabled1562d,
			match=>matchd1562d,
			run=>run);

	Enabled1562d <= matchd1561d;
	-- d1563d
	sted1563d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1563d,
			Enable=>Enabled1563d,
			match=>matchd1563d,
			run=>run);

	Enabled1563d <= matchd1562d OR matchd1563d;
	-- d1564d
	sted1564d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1564d,
			Enable=>Enabled1564d,
			match=>matchd1564d,
			run=>run);

	Enabled1564d <= matchd1563d;
	-- d1565d
	sted1565d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1565d,
			Enable=>Enabled1565d,
			match=>matchd1565d,
			run=>run);

	Enabled1565d <= matchd1564d;
	-- d1566d
	sted1566d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1566d,
			Enable=>Enabled1566d,
			match=>matchd1566d,
			run=>run);

	Enabled1566d <= matchd1565d;
	-- d1567d
	sted1567d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1567d,
			Enable=>Enabled1567d,
			match=>matchd1567d,
			run=>run);

	Enabled1567d <= matchd1566d;
	-- d1568d
	sted1568d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1568d,
			Enable=>Enabled1568d,
			match=>matchd1568d,
			run=>run);

	Enabled1568d <= matchd1567d OR matchd1568d;
	-- d1569d
	sted1569d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1569d,
			Enable=>Enabled1569d,
			match=>matchd1569d,
			run=>run);

	Enabled1569d <= matchd1568d;
	-- d1570d
	sted1570d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1570d,
			Enable=>Enabled1570d,
			match=>matchd1570d,
			run=>run);

	Enabled1570d <= matchd1569d;
	-- d1571d
	sted1571d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1571d,
			Enable=>Enabled1571d,
			match=>matchd1571d,
			run=>run);

	Enabled1571d <= matchd1570d;
	-- d1572d
	sted1572d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1572d,
			Enable=>Enabled1572d,
			match=>matchd1572d,
			run=>run);

	reports(76) <= matchd1572d;
	Enabled1572d <= matchd1571d;
	-- d1573d
	sted1573d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1573d,
			Enable=>Enabled1573d,
			match=>matchd1573d,
			run=>run);

	-- d1574d
	sted1574d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1574d,
			Enable=>Enabled1574d,
			match=>matchd1574d,
			run=>run);

	Enabled1574d <= matchd1573d OR matchd1574d;
	-- d1575d
	sted1575d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1575d,
			Enable=>Enabled1575d,
			match=>matchd1575d,
			run=>run);

	Enabled1575d <= matchd1574d;
	-- d1576d
	sted1576d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1576d,
			Enable=>Enabled1576d,
			match=>matchd1576d,
			run=>run);

	Enabled1576d <= matchd1575d;
	-- d1577d
	sted1577d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1577d,
			Enable=>Enabled1577d,
			match=>matchd1577d,
			run=>run);

	Enabled1577d <= matchd1576d;
	-- d1578d
	sted1578d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1578d,
			Enable=>Enabled1578d,
			match=>matchd1578d,
			run=>run);

	Enabled1578d <= matchd1577d;
	-- d1579d
	sted1579d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1579d,
			Enable=>Enabled1579d,
			match=>matchd1579d,
			run=>run);

	Enabled1579d <= matchd1578d;
	-- d1580d
	sted1580d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1580d,
			Enable=>Enabled1580d,
			match=>matchd1580d,
			run=>run);

	Enabled1580d <= matchd1579d OR matchd1580d;
	-- d1581d
	sted1581d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1581d,
			Enable=>Enabled1581d,
			match=>matchd1581d,
			run=>run);

	Enabled1581d <= matchd1580d;
	-- d1582d
	sted1582d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1582d,
			Enable=>Enabled1582d,
			match=>matchd1582d,
			run=>run);

	Enabled1582d <= matchd1581d;
	-- d1583d
	sted1583d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1583d,
			Enable=>Enabled1583d,
			match=>matchd1583d,
			run=>run);

	Enabled1583d <= matchd1582d;
	-- d1584d
	sted1584d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1584d,
			Enable=>Enabled1584d,
			match=>matchd1584d,
			run=>run);

	reports(77) <= matchd1584d;
	Enabled1584d <= matchd1583d;
	-- d1585d
	sted1585d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1585d,
			Enable=>Enabled1585d,
			match=>matchd1585d,
			run=>run);

	-- d1586d
	sted1586d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1586d,
			Enable=>Enabled1586d,
			match=>matchd1586d,
			run=>run);

	Enabled1586d <= matchd1585d OR matchd1586d;
	-- d1587d
	sted1587d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1587d,
			Enable=>Enabled1587d,
			match=>matchd1587d,
			run=>run);

	Enabled1587d <= matchd1586d;
	-- d1588d
	sted1588d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1588d,
			Enable=>Enabled1588d,
			match=>matchd1588d,
			run=>run);

	Enabled1588d <= matchd1587d;
	-- d1589d
	sted1589d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1589d,
			Enable=>Enabled1589d,
			match=>matchd1589d,
			run=>run);

	Enabled1589d <= matchd1588d;
	-- d1590d
	sted1590d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1590d,
			Enable=>Enabled1590d,
			match=>matchd1590d,
			run=>run);

	Enabled1590d <= matchd1589d;
	-- d1591d
	sted1591d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1591d,
			Enable=>Enabled1591d,
			match=>matchd1591d,
			run=>run);

	Enabled1591d <= matchd1590d;
	-- d1592d
	sted1592d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1592d,
			Enable=>Enabled1592d,
			match=>matchd1592d,
			run=>run);

	Enabled1592d <= matchd1591d;
	-- d1593d
	sted1593d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1593d,
			Enable=>Enabled1593d,
			match=>matchd1593d,
			run=>run);

	Enabled1593d <= matchd1592d;
	-- d1594d
	sted1594d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1594d,
			Enable=>Enabled1594d,
			match=>matchd1594d,
			run=>run);

	Enabled1594d <= matchd1593d;
	-- d1595d
	sted1595d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1595d,
			Enable=>Enabled1595d,
			match=>matchd1595d,
			run=>run);

	Enabled1595d <= matchd1594d;
	-- d1596d
	sted1596d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1596d,
			Enable=>Enabled1596d,
			match=>matchd1596d,
			run=>run);

	Enabled1596d <= matchd1595d;
	-- d1597d
	sted1597d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1597d,
			Enable=>Enabled1597d,
			match=>matchd1597d,
			run=>run);

	Enabled1597d <= matchd1596d;
	-- d1598d
	sted1598d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1598d,
			Enable=>Enabled1598d,
			match=>matchd1598d,
			run=>run);

	reports(78) <= matchd1598d;
	Enabled1598d <= matchd1597d;
	-- d1599d
	sted1599d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1599d,
			Enable=>Enabled1599d,
			match=>matchd1599d,
			run=>run);

	-- d1600d
	sted1600d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1600d,
			Enable=>Enabled1600d,
			match=>matchd1600d,
			run=>run);

	Enabled1600d <= matchd1599d OR matchd1600d;
	-- d1601d
	sted1601d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1601d,
			Enable=>Enabled1601d,
			match=>matchd1601d,
			run=>run);

	Enabled1601d <= matchd1600d;
	-- d1602d
	sted1602d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1602d,
			Enable=>Enabled1602d,
			match=>matchd1602d,
			run=>run);

	Enabled1602d <= matchd1601d;
	-- d1603d
	sted1603d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1603d,
			Enable=>Enabled1603d,
			match=>matchd1603d,
			run=>run);

	Enabled1603d <= matchd1602d;
	-- d1604d
	sted1604d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1604d,
			Enable=>Enabled1604d,
			match=>matchd1604d,
			run=>run);

	Enabled1604d <= matchd1603d;
	-- d1605d
	sted1605d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1605d,
			Enable=>Enabled1605d,
			match=>matchd1605d,
			run=>run);

	Enabled1605d <= matchd1605d OR matchd1604d;
	-- d1606d
	sted1606d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1606d,
			Enable=>Enabled1606d,
			match=>matchd1606d,
			run=>run);

	Enabled1606d <= matchd1605d;
	-- d1607d
	sted1607d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1607d,
			Enable=>Enabled1607d,
			match=>matchd1607d,
			run=>run);

	Enabled1607d <= matchd1606d;
	-- d1608d
	sted1608d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1608d,
			Enable=>Enabled1608d,
			match=>matchd1608d,
			run=>run);

	Enabled1608d <= matchd1607d;
	-- d1609d
	sted1609d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1609d,
			Enable=>Enabled1609d,
			match=>matchd1609d,
			run=>run);

	reports(79) <= matchd1609d;
	Enabled1609d <= matchd1608d;
	-- d1610d
	sted1610d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1610d,
			Enable=>Enabled1610d,
			match=>matchd1610d,
			run=>run);

	-- d1611d
	sted1611d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1611d,
			Enable=>Enabled1611d,
			match=>matchd1611d,
			run=>run);

	Enabled1611d <= matchd1610d OR matchd1611d;
	-- d1612d
	sted1612d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1612d,
			Enable=>Enabled1612d,
			match=>matchd1612d,
			run=>run);

	Enabled1612d <= matchd1611d;
	-- d1613d
	sted1613d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1613d,
			Enable=>Enabled1613d,
			match=>matchd1613d,
			run=>run);

	Enabled1613d <= matchd1612d;
	-- d1614d
	sted1614d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1614d,
			Enable=>Enabled1614d,
			match=>matchd1614d,
			run=>run);

	Enabled1614d <= matchd1613d;
	-- d1615d
	sted1615d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1615d,
			Enable=>Enabled1615d,
			match=>matchd1615d,
			run=>run);

	Enabled1615d <= matchd1614d;
	-- d1616d
	sted1616d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1616d,
			Enable=>Enabled1616d,
			match=>matchd1616d,
			run=>run);

	Enabled1616d <= matchd1615d;
	-- d1617d
	sted1617d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1617d,
			Enable=>Enabled1617d,
			match=>matchd1617d,
			run=>run);

	Enabled1617d <= matchd1617d OR matchd1616d;
	-- d1618d
	sted1618d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1618d,
			Enable=>Enabled1618d,
			match=>matchd1618d,
			run=>run);

	Enabled1618d <= matchd1617d;
	-- d1619d
	sted1619d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1619d,
			Enable=>Enabled1619d,
			match=>matchd1619d,
			run=>run);

	Enabled1619d <= matchd1618d;
	-- d1620d
	sted1620d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1620d,
			Enable=>Enabled1620d,
			match=>matchd1620d,
			run=>run);

	Enabled1620d <= matchd1619d;
	-- d1621d
	sted1621d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1621d,
			Enable=>Enabled1621d,
			match=>matchd1621d,
			run=>run);

	reports(80) <= matchd1621d;
	Enabled1621d <= matchd1620d;
	-- d1622d
	sted1622d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1622d,
			Enable=>Enabled1622d,
			match=>matchd1622d,
			run=>run);

	-- d1623d
	sted1623d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1623d,
			Enable=>Enabled1623d,
			match=>matchd1623d,
			run=>run);

	Enabled1623d <= matchd1622d;
	-- d1624d
	sted1624d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1624d,
			Enable=>Enabled1624d,
			match=>matchd1624d,
			run=>run);

	Enabled1624d <= matchd1623d;
	-- d1625d
	sted1625d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1625d,
			Enable=>Enabled1625d,
			match=>matchd1625d,
			run=>run);

	Enabled1625d <= matchd1624d;
	-- d1626d
	sted1626d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1626d,
			Enable=>Enabled1626d,
			match=>matchd1626d,
			run=>run);

	Enabled1626d <= matchd1625d;
	-- d1627d
	sted1627d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1627d,
			Enable=>Enabled1627d,
			match=>matchd1627d,
			run=>run);

	Enabled1627d <= matchd1626d;
	-- d1628d
	sted1628d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1628d,
			Enable=>Enabled1628d,
			match=>matchd1628d,
			run=>run);

	Enabled1628d <= matchd1627d;
	-- d1629d
	sted1629d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1629d,
			Enable=>Enabled1629d,
			match=>matchd1629d,
			run=>run);

	Enabled1629d <= matchd1628d;
	-- d1630d
	sted1630d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1630d,
			Enable=>Enabled1630d,
			match=>matchd1630d,
			run=>run);

	reports(81) <= matchd1630d;
	Enabled1630d <= matchd1629d;
	-- d1631d
	sted1631d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1631d,
			Enable=>Enabled1631d,
			match=>matchd1631d,
			run=>run);

	-- d1632d
	sted1632d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1632d,
			Enable=>Enabled1632d,
			match=>matchd1632d,
			run=>run);

	Enabled1632d <= matchd1631d OR matchd1632d;
	-- d1633d
	sted1633d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1633d,
			Enable=>Enabled1633d,
			match=>matchd1633d,
			run=>run);

	Enabled1633d <= matchd1632d;
	-- d1634d
	sted1634d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1634d,
			Enable=>Enabled1634d,
			match=>matchd1634d,
			run=>run);

	Enabled1634d <= matchd1633d;
	-- d1635d
	sted1635d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1635d,
			Enable=>Enabled1635d,
			match=>matchd1635d,
			run=>run);

	Enabled1635d <= matchd1634d;
	-- d1636d
	sted1636d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1636d,
			Enable=>Enabled1636d,
			match=>matchd1636d,
			run=>run);

	Enabled1636d <= matchd1635d;
	-- d1637d
	sted1637d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1637d,
			Enable=>Enabled1637d,
			match=>matchd1637d,
			run=>run);

	Enabled1637d <= matchd1636d OR matchd1637d;
	-- d1638d
	sted1638d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1638d,
			Enable=>Enabled1638d,
			match=>matchd1638d,
			run=>run);

	Enabled1638d <= matchd1637d;
	-- d1639d
	sted1639d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1639d,
			Enable=>Enabled1639d,
			match=>matchd1639d,
			run=>run);

	Enabled1639d <= matchd1638d;
	-- d1640d
	sted1640d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1640d,
			Enable=>Enabled1640d,
			match=>matchd1640d,
			run=>run);

	Enabled1640d <= matchd1639d;
	-- d1641d
	sted1641d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1641d,
			Enable=>Enabled1641d,
			match=>matchd1641d,
			run=>run);

	Enabled1641d <= matchd1640d;
	-- d1642d
	sted1642d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1642d,
			Enable=>Enabled1642d,
			match=>matchd1642d,
			run=>run);

	reports(82) <= matchd1642d;
	Enabled1642d <= matchd1641d;
	-- d1643d
	sted1643d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1643d,
			Enable=>Enabled1643d,
			match=>matchd1643d,
			run=>run);

	-- d1644d
	sted1644d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1644d,
			Enable=>Enabled1644d,
			match=>matchd1644d,
			run=>run);

	Enabled1644d <= matchd1644d OR matchd1643d;
	-- d1645d
	sted1645d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1645d,
			Enable=>Enabled1645d,
			match=>matchd1645d,
			run=>run);

	Enabled1645d <= matchd1644d;
	-- d1646d
	sted1646d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1646d,
			Enable=>Enabled1646d,
			match=>matchd1646d,
			run=>run);

	Enabled1646d <= matchd1645d;
	-- d1647d
	sted1647d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1647d,
			Enable=>Enabled1647d,
			match=>matchd1647d,
			run=>run);

	Enabled1647d <= matchd1646d;
	-- d1648d
	sted1648d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1648d,
			Enable=>Enabled1648d,
			match=>matchd1648d,
			run=>run);

	Enabled1648d <= matchd1647d;
	-- d1649d
	sted1649d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1649d,
			Enable=>Enabled1649d,
			match=>matchd1649d,
			run=>run);

	Enabled1649d <= matchd1649d OR matchd1648d;
	-- d1650d
	sted1650d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1650d,
			Enable=>Enabled1650d,
			match=>matchd1650d,
			run=>run);

	Enabled1650d <= matchd1649d;
	-- d1651d
	sted1651d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1651d,
			Enable=>Enabled1651d,
			match=>matchd1651d,
			run=>run);

	Enabled1651d <= matchd1650d;
	-- d1652d
	sted1652d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1652d,
			Enable=>Enabled1652d,
			match=>matchd1652d,
			run=>run);

	Enabled1652d <= matchd1651d;
	-- d1653d
	sted1653d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1653d,
			Enable=>Enabled1653d,
			match=>matchd1653d,
			run=>run);

	reports(83) <= matchd1653d;
	Enabled1653d <= matchd1652d;
	-- d1654d
	sted1654d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1654d,
			Enable=>Enabled1654d,
			match=>matchd1654d,
			run=>run);

	-- d1655d
	sted1655d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1655d,
			Enable=>Enabled1655d,
			match=>matchd1655d,
			run=>run);

	Enabled1655d <= matchd1655d OR matchd1654d;
	-- d1656d
	sted1656d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1656d,
			Enable=>Enabled1656d,
			match=>matchd1656d,
			run=>run);

	Enabled1656d <= matchd1655d;
	-- d1657d
	sted1657d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1657d,
			Enable=>Enabled1657d,
			match=>matchd1657d,
			run=>run);

	Enabled1657d <= matchd1656d;
	-- d1658d
	sted1658d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1658d,
			Enable=>Enabled1658d,
			match=>matchd1658d,
			run=>run);

	Enabled1658d <= matchd1657d;
	-- d1659d
	sted1659d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1659d,
			Enable=>Enabled1659d,
			match=>matchd1659d,
			run=>run);

	Enabled1659d <= matchd1658d;
	-- d1660d
	sted1660d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1660d,
			Enable=>Enabled1660d,
			match=>matchd1660d,
			run=>run);

	Enabled1660d <= matchd1659d;
	-- d1661d
	sted1661d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1661d,
			Enable=>Enabled1661d,
			match=>matchd1661d,
			run=>run);

	Enabled1661d <= matchd1660d;
	-- d1662d
	sted1662d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1662d,
			Enable=>Enabled1662d,
			match=>matchd1662d,
			run=>run);

	Enabled1662d <= matchd1661d;
	-- d1663d
	sted1663d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1663d,
			Enable=>Enabled1663d,
			match=>matchd1663d,
			run=>run);

	Enabled1663d <= matchd1662d;
	-- d1664d
	sted1664d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1664d,
			Enable=>Enabled1664d,
			match=>matchd1664d,
			run=>run);

	Enabled1664d <= matchd1664d OR matchd1663d;
	-- d1665d
	sted1665d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1665d,
			Enable=>Enabled1665d,
			match=>matchd1665d,
			run=>run);

	Enabled1665d <= matchd1664d;
	-- d1666d
	sted1666d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1666d,
			Enable=>Enabled1666d,
			match=>matchd1666d,
			run=>run);

	Enabled1666d <= matchd1665d;
	-- d1667d
	sted1667d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1667d,
			Enable=>Enabled1667d,
			match=>matchd1667d,
			run=>run);

	Enabled1667d <= matchd1666d;
	-- d1668d
	sted1668d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1668d,
			Enable=>Enabled1668d,
			match=>matchd1668d,
			run=>run);

	Enabled1668d <= matchd1667d;
	-- d1669d
	sted1669d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1669d,
			Enable=>Enabled1669d,
			match=>matchd1669d,
			run=>run);

	Enabled1669d <= matchd1669d OR matchd1668d;
	-- d1670d
	sted1670d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1670d,
			Enable=>Enabled1670d,
			match=>matchd1670d,
			run=>run);

	Enabled1670d <= matchd1669d;
	-- d1671d
	sted1671d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1671d,
			Enable=>Enabled1671d,
			match=>matchd1671d,
			run=>run);

	Enabled1671d <= matchd1670d;
	-- d1672d
	sted1672d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1672d,
			Enable=>Enabled1672d,
			match=>matchd1672d,
			run=>run);

	reports(84) <= matchd1672d;
	Enabled1672d <= matchd1671d;
	-- d1673d
	sted1673d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1673d,
			Enable=>Enabled1673d,
			match=>matchd1673d,
			run=>run);

	-- d1674d
	sted1674d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1674d,
			Enable=>Enabled1674d,
			match=>matchd1674d,
			run=>run);

	Enabled1674d <= matchd1673d OR matchd1674d;
	-- d1675d
	sted1675d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1675d,
			Enable=>Enabled1675d,
			match=>matchd1675d,
			run=>run);

	Enabled1675d <= matchd1674d;
	-- d1676d
	sted1676d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1676d,
			Enable=>Enabled1676d,
			match=>matchd1676d,
			run=>run);

	Enabled1676d <= matchd1675d;
	-- d1677d
	sted1677d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1677d,
			Enable=>Enabled1677d,
			match=>matchd1677d,
			run=>run);

	Enabled1677d <= matchd1676d;
	-- d1678d
	sted1678d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1678d,
			Enable=>Enabled1678d,
			match=>matchd1678d,
			run=>run);

	Enabled1678d <= matchd1677d;
	-- d1679d
	sted1679d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1679d,
			Enable=>Enabled1679d,
			match=>matchd1679d,
			run=>run);

	Enabled1679d <= matchd1678d OR matchd1679d;
	-- d1680d
	sted1680d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1680d,
			Enable=>Enabled1680d,
			match=>matchd1680d,
			run=>run);

	Enabled1680d <= matchd1679d;
	-- d1681d
	sted1681d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1681d,
			Enable=>Enabled1681d,
			match=>matchd1681d,
			run=>run);

	Enabled1681d <= matchd1680d;
	-- d1682d
	sted1682d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1682d,
			Enable=>Enabled1682d,
			match=>matchd1682d,
			run=>run);

	Enabled1682d <= matchd1681d;
	-- d1683d
	sted1683d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1683d,
			Enable=>Enabled1683d,
			match=>matchd1683d,
			run=>run);

	Enabled1683d <= matchd1682d;
	-- d1684d
	sted1684d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1684d,
			Enable=>Enabled1684d,
			match=>matchd1684d,
			run=>run);

	Enabled1684d <= matchd1683d;
	-- d1685d
	sted1685d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1685d,
			Enable=>Enabled1685d,
			match=>matchd1685d,
			run=>run);

	Enabled1685d <= matchd1684d OR matchd1685d;
	-- d1686d
	sted1686d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1686d,
			Enable=>Enabled1686d,
			match=>matchd1686d,
			run=>run);

	Enabled1686d <= matchd1685d;
	-- d1687d
	sted1687d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1687d,
			Enable=>Enabled1687d,
			match=>matchd1687d,
			run=>run);

	Enabled1687d <= matchd1686d;
	-- d1688d
	sted1688d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1688d,
			Enable=>Enabled1688d,
			match=>matchd1688d,
			run=>run);

	Enabled1688d <= matchd1687d;
	-- d1689d
	sted1689d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1689d,
			Enable=>Enabled1689d,
			match=>matchd1689d,
			run=>run);

	Enabled1689d <= matchd1688d;
	-- d1690d
	sted1690d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1690d,
			Enable=>Enabled1690d,
			match=>matchd1690d,
			run=>run);

	reports(85) <= matchd1690d;
	Enabled1690d <= matchd1689d;
	-- d1691d
	sted1691d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1691d,
			Enable=>Enabled1691d,
			match=>matchd1691d,
			run=>run);

	-- d1692d
	sted1692d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1692d,
			Enable=>Enabled1692d,
			match=>matchd1692d,
			run=>run);

	Enabled1692d <= matchd1692d OR matchd1691d;
	-- d1693d
	sted1693d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1693d,
			Enable=>Enabled1693d,
			match=>matchd1693d,
			run=>run);

	Enabled1693d <= matchd1692d;
	-- d1694d
	sted1694d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1694d,
			Enable=>Enabled1694d,
			match=>matchd1694d,
			run=>run);

	Enabled1694d <= matchd1693d;
	-- d1695d
	sted1695d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1695d,
			Enable=>Enabled1695d,
			match=>matchd1695d,
			run=>run);

	Enabled1695d <= matchd1694d;
	-- d1696d
	sted1696d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1696d,
			Enable=>Enabled1696d,
			match=>matchd1696d,
			run=>run);

	Enabled1696d <= matchd1695d;
	-- d1697d
	sted1697d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1697d,
			Enable=>Enabled1697d,
			match=>matchd1697d,
			run=>run);

	Enabled1697d <= matchd1697d OR matchd1696d;
	-- d1698d
	sted1698d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1698d,
			Enable=>Enabled1698d,
			match=>matchd1698d,
			run=>run);

	Enabled1698d <= matchd1697d;
	-- d1699d
	sted1699d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1699d,
			Enable=>Enabled1699d,
			match=>matchd1699d,
			run=>run);

	Enabled1699d <= matchd1698d;
	-- d1700d
	sted1700d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1700d,
			Enable=>Enabled1700d,
			match=>matchd1700d,
			run=>run);

	Enabled1700d <= matchd1699d;
	-- d1701d
	sted1701d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1701d,
			Enable=>Enabled1701d,
			match=>matchd1701d,
			run=>run);

	reports(86) <= matchd1701d;
	Enabled1701d <= matchd1700d;
	-- d1702d
	sted1702d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1702d,
			Enable=>Enabled1702d,
			match=>matchd1702d,
			run=>run);

	-- d1703d
	sted1703d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1703d,
			Enable=>Enabled1703d,
			match=>matchd1703d,
			run=>run);

	Enabled1703d <= matchd1702d OR matchd1703d;
	-- d1704d
	sted1704d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1704d,
			Enable=>Enabled1704d,
			match=>matchd1704d,
			run=>run);

	Enabled1704d <= matchd1703d;
	-- d1705d
	sted1705d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1705d,
			Enable=>Enabled1705d,
			match=>matchd1705d,
			run=>run);

	Enabled1705d <= matchd1704d;
	-- d1706d
	sted1706d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1706d,
			Enable=>Enabled1706d,
			match=>matchd1706d,
			run=>run);

	Enabled1706d <= matchd1705d;
	-- d1707d
	sted1707d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1707d,
			Enable=>Enabled1707d,
			match=>matchd1707d,
			run=>run);

	Enabled1707d <= matchd1706d;
	-- d1708d
	sted1708d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1708d,
			Enable=>Enabled1708d,
			match=>matchd1708d,
			run=>run);

	Enabled1708d <= matchd1707d OR matchd1708d;
	-- d1709d
	sted1709d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1709d,
			Enable=>Enabled1709d,
			match=>matchd1709d,
			run=>run);

	Enabled1709d <= matchd1708d;
	-- d1710d
	sted1710d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1710d,
			Enable=>Enabled1710d,
			match=>matchd1710d,
			run=>run);

	Enabled1710d <= matchd1709d;
	-- d1711d
	sted1711d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1711d,
			Enable=>Enabled1711d,
			match=>matchd1711d,
			run=>run);

	Enabled1711d <= matchd1710d;
	-- d1712d
	sted1712d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1712d,
			Enable=>Enabled1712d,
			match=>matchd1712d,
			run=>run);

	Enabled1712d <= matchd1711d;
	-- d1713d
	sted1713d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1713d,
			Enable=>Enabled1713d,
			match=>matchd1713d,
			run=>run);

	Enabled1713d <= matchd1713d OR matchd1712d;
	-- d1714d
	sted1714d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1714d,
			Enable=>Enabled1714d,
			match=>matchd1714d,
			run=>run);

	Enabled1714d <= matchd1713d;
	-- d1715d
	sted1715d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1715d,
			Enable=>Enabled1715d,
			match=>matchd1715d,
			run=>run);

	Enabled1715d <= matchd1714d;
	-- d1716d
	sted1716d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1716d,
			Enable=>Enabled1716d,
			match=>matchd1716d,
			run=>run);

	reports(87) <= matchd1716d;
	Enabled1716d <= matchd1715d;
	-- d1717d
	sted1717d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1717d,
			Enable=>Enabled1717d,
			match=>matchd1717d,
			run=>run);

	-- d1718d
	sted1718d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1718d,
			Enable=>Enabled1718d,
			match=>matchd1718d,
			run=>run);

	Enabled1718d <= matchd1717d OR matchd1718d;
	-- d1719d
	sted1719d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1719d,
			Enable=>Enabled1719d,
			match=>matchd1719d,
			run=>run);

	Enabled1719d <= matchd1718d;
	-- d1720d
	sted1720d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1720d,
			Enable=>Enabled1720d,
			match=>matchd1720d,
			run=>run);

	Enabled1720d <= matchd1719d;
	-- d1721d
	sted1721d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1721d,
			Enable=>Enabled1721d,
			match=>matchd1721d,
			run=>run);

	Enabled1721d <= matchd1720d;
	-- d1722d
	sted1722d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1722d,
			Enable=>Enabled1722d,
			match=>matchd1722d,
			run=>run);

	Enabled1722d <= matchd1721d;
	-- d1723d
	sted1723d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1723d,
			Enable=>Enabled1723d,
			match=>matchd1723d,
			run=>run);

	Enabled1723d <= matchd1722d OR matchd1723d;
	-- d1724d
	sted1724d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1724d,
			Enable=>Enabled1724d,
			match=>matchd1724d,
			run=>run);

	Enabled1724d <= matchd1723d;
	-- d1725d
	sted1725d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1725d,
			Enable=>Enabled1725d,
			match=>matchd1725d,
			run=>run);

	Enabled1725d <= matchd1724d;
	-- d1726d
	sted1726d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1726d,
			Enable=>Enabled1726d,
			match=>matchd1726d,
			run=>run);

	Enabled1726d <= matchd1725d;
	-- d1727d
	sted1727d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1727d,
			Enable=>Enabled1727d,
			match=>matchd1727d,
			run=>run);

	Enabled1727d <= matchd1726d;
	-- d1728d
	sted1728d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1728d,
			Enable=>Enabled1728d,
			match=>matchd1728d,
			run=>run);

	reports(88) <= matchd1728d;
	Enabled1728d <= matchd1727d;
	-- d1729d
	sted1729d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1729d,
			Enable=>Enabled1729d,
			match=>matchd1729d,
			run=>run);

	-- d1730d
	sted1730d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1730d,
			Enable=>Enabled1730d,
			match=>matchd1730d,
			run=>run);

	Enabled1730d <= matchd1729d OR matchd1730d;
	-- d1731d
	sted1731d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1731d,
			Enable=>Enabled1731d,
			match=>matchd1731d,
			run=>run);

	Enabled1731d <= matchd1730d;
	-- d1732d
	sted1732d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1732d,
			Enable=>Enabled1732d,
			match=>matchd1732d,
			run=>run);

	Enabled1732d <= matchd1731d OR matchd1732d;
	-- d1733d
	sted1733d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1733d,
			Enable=>Enabled1733d,
			match=>matchd1733d,
			run=>run);

	Enabled1733d <= matchd1732d;
	-- d1734d
	sted1734d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1734d,
			Enable=>Enabled1734d,
			match=>matchd1734d,
			run=>run);

	Enabled1734d <= matchd1733d;
	-- d1735d
	sted1735d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1735d,
			Enable=>Enabled1735d,
			match=>matchd1735d,
			run=>run);

	Enabled1735d <= matchd1734d;
	-- d1736d
	sted1736d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1736d,
			Enable=>Enabled1736d,
			match=>matchd1736d,
			run=>run);

	Enabled1736d <= matchd1735d;
	-- d1737d
	sted1737d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1737d,
			Enable=>Enabled1737d,
			match=>matchd1737d,
			run=>run);

	Enabled1737d <= matchd1736d;
	-- d1738d
	sted1738d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1738d,
			Enable=>Enabled1738d,
			match=>matchd1738d,
			run=>run);

	Enabled1738d <= matchd1737d;
	-- d1739d
	sted1739d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1739d,
			Enable=>Enabled1739d,
			match=>matchd1739d,
			run=>run);

	Enabled1739d <= matchd1739d OR matchd1738d;
	-- d1740d
	sted1740d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1740d,
			Enable=>Enabled1740d,
			match=>matchd1740d,
			run=>run);

	Enabled1740d <= matchd1739d;
	-- d1741d
	sted1741d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1741d,
			Enable=>Enabled1741d,
			match=>matchd1741d,
			run=>run);

	Enabled1741d <= matchd1740d OR matchd1741d;
	-- d1742d
	sted1742d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1742d,
			Enable=>Enabled1742d,
			match=>matchd1742d,
			run=>run);

	Enabled1742d <= matchd1741d;
	-- d1743d
	sted1743d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1743d,
			Enable=>Enabled1743d,
			match=>matchd1743d,
			run=>run);

	Enabled1743d <= matchd1742d;
	-- d1744d
	sted1744d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1744d,
			Enable=>Enabled1744d,
			match=>matchd1744d,
			run=>run);

	Enabled1744d <= matchd1743d;
	-- d1745d
	sted1745d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1745d,
			Enable=>Enabled1745d,
			match=>matchd1745d,
			run=>run);

	Enabled1745d <= matchd1744d;
	-- d1746d
	sted1746d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1746d,
			Enable=>Enabled1746d,
			match=>matchd1746d,
			run=>run);

	-- d1747d
	sted1747d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1747d,
			Enable=>Enabled1747d,
			match=>matchd1747d,
			run=>run);

	Enabled1747d <= matchd1746d;
	-- d1748d
	sted1748d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1748d,
			Enable=>Enabled1748d,
			match=>matchd1748d,
			run=>run);

	Enabled1748d <= matchd1747d;
	-- d1749d
	sted1749d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1749d,
			Enable=>Enabled1749d,
			match=>matchd1749d,
			run=>run);

	Enabled1749d <= matchd1748d;
	-- d1750d
	sted1750d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1750d,
			Enable=>Enabled1750d,
			match=>matchd1750d,
			run=>run);

	Enabled1750d <= matchd1749d;
	-- d1751d
	sted1751d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1751d,
			Enable=>Enabled1751d,
			match=>matchd1751d,
			run=>run);

	Enabled1751d <= matchd1750d;
	-- d1752d
	sted1752d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1752d,
			Enable=>Enabled1752d,
			match=>matchd1752d,
			run=>run);

	Enabled1752d <= matchd1752d OR matchd1751d;
	-- d1753d
	sted1753d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1753d,
			Enable=>Enabled1753d,
			match=>matchd1753d,
			run=>run);

	Enabled1753d <= matchd1752d;
	-- d1754d
	sted1754d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1754d,
			Enable=>Enabled1754d,
			match=>matchd1754d,
			run=>run);

	Enabled1754d <= matchd1754d OR matchd1753d;
	-- d1755d
	sted1755d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1755d,
			Enable=>Enabled1755d,
			match=>matchd1755d,
			run=>run);

	Enabled1755d <= matchd1754d;
	-- d1756d
	sted1756d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1756d,
			Enable=>Enabled1756d,
			match=>matchd1756d,
			run=>run);

	Enabled1756d <= matchd1756d OR matchd1755d;
	-- d1757d
	sted1757d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1757d,
			Enable=>Enabled1757d,
			match=>matchd1757d,
			run=>run);

	Enabled1757d <= matchd1756d;
	-- d1758d
	sted1758d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1758d,
			Enable=>Enabled1758d,
			match=>matchd1758d,
			run=>run);

	Enabled1758d <= matchd1758d OR matchd1757d;
	-- d1759d
	sted1759d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1759d,
			Enable=>Enabled1759d,
			match=>matchd1759d,
			run=>run);

	Enabled1759d <= matchd1758d;
	-- d1760d
	sted1760d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1760d,
			Enable=>Enabled1760d,
			match=>matchd1760d,
			run=>run);

	Enabled1760d <= matchd1759d;
	-- d1761d
	sted1761d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1761d,
			Enable=>Enabled1761d,
			match=>matchd1761d,
			run=>run);

	Enabled1761d <= matchd1760d;
	-- d1762d
	sted1762d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1762d,
			Enable=>Enabled1762d,
			match=>matchd1762d,
			run=>run);

	Enabled1762d <= matchd1761d;
	-- d1764d
	sted1764d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1764d,
			Enable=>Enabled1764d,
			match=>matchd1764d,
			run=>run);

	-- d1765d
	sted1765d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1765d,
			Enable=>Enabled1765d,
			match=>matchd1765d,
			run=>run);

	Enabled1765d <= matchd1764d OR matchd1765d;
	-- d1766d
	sted1766d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1766d,
			Enable=>Enabled1766d,
			match=>matchd1766d,
			run=>run);

	Enabled1766d <= matchd1765d;
	-- d1767d
	sted1767d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1767d,
			Enable=>Enabled1767d,
			match=>matchd1767d,
			run=>run);

	Enabled1767d <= matchd1766d;
	-- d1768d
	sted1768d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1768d,
			Enable=>Enabled1768d,
			match=>matchd1768d,
			run=>run);

	Enabled1768d <= matchd1767d;
	-- d1769d
	sted1769d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1769d,
			Enable=>Enabled1769d,
			match=>matchd1769d,
			run=>run);

	Enabled1769d <= matchd1768d;
	-- d1770d
	sted1770d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1770d,
			Enable=>Enabled1770d,
			match=>matchd1770d,
			run=>run);

	Enabled1770d <= matchd1769d OR matchd1770d;
	-- d1771d
	sted1771d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1771d,
			Enable=>Enabled1771d,
			match=>matchd1771d,
			run=>run);

	Enabled1771d <= matchd1770d;
	-- d1772d
	sted1772d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1772d,
			Enable=>Enabled1772d,
			match=>matchd1772d,
			run=>run);

	Enabled1772d <= matchd1771d;
	-- d1773d
	sted1773d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1773d,
			Enable=>Enabled1773d,
			match=>matchd1773d,
			run=>run);

	Enabled1773d <= matchd1772d;
	-- d1774d
	sted1774d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1774d,
			Enable=>Enabled1774d,
			match=>matchd1774d,
			run=>run);

	reports(89) <= matchd1774d;
	Enabled1774d <= matchd1773d;
	-- d1775d
	sted1775d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1775d,
			Enable=>Enabled1775d,
			match=>matchd1775d,
			run=>run);

	-- d1776d
	sted1776d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1776d,
			Enable=>Enabled1776d,
			match=>matchd1776d,
			run=>run);

	Enabled1776d <= matchd1776d OR matchd1775d;
	-- d1777d
	sted1777d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1777d,
			Enable=>Enabled1777d,
			match=>matchd1777d,
			run=>run);

	Enabled1777d <= matchd1776d;
	-- d1778d
	sted1778d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1778d,
			Enable=>Enabled1778d,
			match=>matchd1778d,
			run=>run);

	Enabled1778d <= matchd1777d;
	-- d1779d
	sted1779d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1779d,
			Enable=>Enabled1779d,
			match=>matchd1779d,
			run=>run);

	Enabled1779d <= matchd1778d;
	-- d1780d
	sted1780d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1780d,
			Enable=>Enabled1780d,
			match=>matchd1780d,
			run=>run);

	Enabled1780d <= matchd1779d;
	-- d1781d
	sted1781d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1781d,
			Enable=>Enabled1781d,
			match=>matchd1781d,
			run=>run);

	Enabled1781d <= matchd1780d;
	-- d1782d
	sted1782d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1782d,
			Enable=>Enabled1782d,
			match=>matchd1782d,
			run=>run);

	Enabled1782d <= matchd1781d;
	-- d1783d
	sted1783d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1783d,
			Enable=>Enabled1783d,
			match=>matchd1783d,
			run=>run);

	Enabled1783d <= matchd1782d;
	-- d1784d
	sted1784d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1784d,
			Enable=>Enabled1784d,
			match=>matchd1784d,
			run=>run);

	Enabled1784d <= matchd1783d OR matchd1784d;
	-- d1785d
	sted1785d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1785d,
			Enable=>Enabled1785d,
			match=>matchd1785d,
			run=>run);

	Enabled1785d <= matchd1784d;
	-- d1786d
	sted1786d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1786d,
			Enable=>Enabled1786d,
			match=>matchd1786d,
			run=>run);

	Enabled1786d <= matchd1785d;
	-- d1787d
	sted1787d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1787d,
			Enable=>Enabled1787d,
			match=>matchd1787d,
			run=>run);

	Enabled1787d <= matchd1786d;
	-- d1788d
	sted1788d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1788d,
			Enable=>Enabled1788d,
			match=>matchd1788d,
			run=>run);

	Enabled1788d <= matchd1787d;
	-- d1789d
	sted1789d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1789d,
			Enable=>Enabled1789d,
			match=>matchd1789d,
			run=>run);

	Enabled1789d <= matchd1788d OR matchd1789d;
	-- d1790d
	sted1790d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1790d,
			Enable=>Enabled1790d,
			match=>matchd1790d,
			run=>run);

	Enabled1790d <= matchd1789d;
	-- d1791d
	sted1791d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1791d,
			Enable=>Enabled1791d,
			match=>matchd1791d,
			run=>run);

	Enabled1791d <= matchd1790d;
	-- d1792d
	sted1792d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1792d,
			Enable=>Enabled1792d,
			match=>matchd1792d,
			run=>run);

	Enabled1792d <= matchd1791d;
	-- d1793d
	sted1793d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1793d,
			Enable=>Enabled1793d,
			match=>matchd1793d,
			run=>run);

	Enabled1793d <= matchd1792d;
	-- d1794d
	sted1794d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1794d,
			Enable=>Enabled1794d,
			match=>matchd1794d,
			run=>run);

	Enabled1794d <= matchd1793d;
	-- d1795d
	sted1795d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1795d,
			Enable=>Enabled1795d,
			match=>matchd1795d,
			run=>run);

	Enabled1795d <= matchd1794d;
	-- d1796d
	sted1796d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1796d,
			Enable=>Enabled1796d,
			match=>matchd1796d,
			run=>run);

	reports(90) <= matchd1796d;
	Enabled1796d <= matchd1795d;
	-- d1797d
	sted1797d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1797d,
			Enable=>Enabled1797d,
			match=>matchd1797d,
			run=>run);

	-- d1798d
	sted1798d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1798d,
			Enable=>Enabled1798d,
			match=>matchd1798d,
			run=>run);

	Enabled1798d <= matchd1797d OR matchd1798d;
	-- d1799d
	sted1799d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1799d,
			Enable=>Enabled1799d,
			match=>matchd1799d,
			run=>run);

	Enabled1799d <= matchd1798d;
	-- d1800d
	sted1800d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1800d,
			Enable=>Enabled1800d,
			match=>matchd1800d,
			run=>run);

	Enabled1800d <= matchd1799d;
	-- d1801d
	sted1801d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1801d,
			Enable=>Enabled1801d,
			match=>matchd1801d,
			run=>run);

	Enabled1801d <= matchd1800d;
	-- d1802d
	sted1802d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1802d,
			Enable=>Enabled1802d,
			match=>matchd1802d,
			run=>run);

	Enabled1802d <= matchd1801d;
	-- d1803d
	sted1803d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1803d,
			Enable=>Enabled1803d,
			match=>matchd1803d,
			run=>run);

	Enabled1803d <= matchd1802d OR matchd1803d;
	-- d1804d
	sted1804d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1804d,
			Enable=>Enabled1804d,
			match=>matchd1804d,
			run=>run);

	Enabled1804d <= matchd1803d;
	-- d1805d
	sted1805d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1805d,
			Enable=>Enabled1805d,
			match=>matchd1805d,
			run=>run);

	Enabled1805d <= matchd1804d;
	-- d1806d
	sted1806d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1806d,
			Enable=>Enabled1806d,
			match=>matchd1806d,
			run=>run);

	Enabled1806d <= matchd1805d;
	-- d1807d
	sted1807d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1807d,
			Enable=>Enabled1807d,
			match=>matchd1807d,
			run=>run);

	Enabled1807d <= matchd1807d OR matchd1806d;
	-- d1808d
	sted1808d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1808d,
			Enable=>Enabled1808d,
			match=>matchd1808d,
			run=>run);

	Enabled1808d <= matchd1807d;
	-- d1809d
	sted1809d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1809d,
			Enable=>Enabled1809d,
			match=>matchd1809d,
			run=>run);

	Enabled1809d <= matchd1809d OR matchd1808d;
	-- d1810d
	sted1810d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1810d,
			Enable=>Enabled1810d,
			match=>matchd1810d,
			run=>run);

	Enabled1810d <= matchd1809d;
	-- d1811d
	sted1811d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1811d,
			Enable=>Enabled1811d,
			match=>matchd1811d,
			run=>run);

	Enabled1811d <= matchd1810d OR matchd1811d;
	-- d1812d
	sted1812d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1812d,
			Enable=>Enabled1812d,
			match=>matchd1812d,
			run=>run);

	Enabled1812d <= matchd1811d;
	-- d1813d
	sted1813d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1813d,
			Enable=>Enabled1813d,
			match=>matchd1813d,
			run=>run);

	Enabled1813d <= matchd1812d OR matchd1813d;
	-- d1814d
	sted1814d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1814d,
			Enable=>Enabled1814d,
			match=>matchd1814d,
			run=>run);

	Enabled1814d <= matchd1813d;
	-- d1815d
	sted1815d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1815d,
			Enable=>Enabled1815d,
			match=>matchd1815d,
			run=>run);

	-- d1816d
	sted1816d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1816d,
			Enable=>Enabled1816d,
			match=>matchd1816d,
			run=>run);

	Enabled1816d <= matchd1816d OR matchd1815d;
	-- d1817d
	sted1817d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1817d,
			Enable=>Enabled1817d,
			match=>matchd1817d,
			run=>run);

	Enabled1817d <= matchd1816d;
	-- d1818d
	sted1818d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1818d,
			Enable=>Enabled1818d,
			match=>matchd1818d,
			run=>run);

	Enabled1818d <= matchd1817d;
	-- d1819d
	sted1819d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1819d,
			Enable=>Enabled1819d,
			match=>matchd1819d,
			run=>run);

	Enabled1819d <= matchd1818d;
	-- d1820d
	sted1820d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1820d,
			Enable=>Enabled1820d,
			match=>matchd1820d,
			run=>run);

	Enabled1820d <= matchd1819d;
	-- d1821d
	sted1821d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1821d,
			Enable=>Enabled1821d,
			match=>matchd1821d,
			run=>run);

	Enabled1821d <= matchd1820d OR matchd1821d;
	-- d1822d
	sted1822d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1822d,
			Enable=>Enabled1822d,
			match=>matchd1822d,
			run=>run);

	Enabled1822d <= matchd1821d;
	-- d1823d
	sted1823d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1823d,
			Enable=>Enabled1823d,
			match=>matchd1823d,
			run=>run);

	Enabled1823d <= matchd1823d OR matchd1822d;
	-- d1824d
	sted1824d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1824d,
			Enable=>Enabled1824d,
			match=>matchd1824d,
			run=>run);

	Enabled1824d <= matchd1823d;
	-- d1825d
	sted1825d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1825d,
			Enable=>Enabled1825d,
			match=>matchd1825d,
			run=>run);

	Enabled1825d <= matchd1825d OR matchd1824d;
	-- d1826d
	sted1826d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1826d,
			Enable=>Enabled1826d,
			match=>matchd1826d,
			run=>run);

	Enabled1826d <= matchd1825d;
	-- d1827d
	sted1827d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1827d,
			Enable=>Enabled1827d,
			match=>matchd1827d,
			run=>run);

	Enabled1827d <= matchd1826d;
	-- d1828d
	sted1828d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1828d,
			Enable=>Enabled1828d,
			match=>matchd1828d,
			run=>run);

	Enabled1828d <= matchd1827d;
	-- d1829d
	sted1829d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1829d,
			Enable=>Enabled1829d,
			match=>matchd1829d,
			run=>run);

	Enabled1829d <= matchd1829d OR matchd1828d;
	-- d1830d
	sted1830d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1830d,
			Enable=>Enabled1830d,
			match=>matchd1830d,
			run=>run);

	Enabled1830d <= matchd1829d;
	-- d1831d
	sted1831d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1831d,
			Enable=>Enabled1831d,
			match=>matchd1831d,
			run=>run);

	Enabled1831d <= matchd1831d OR matchd1830d;
	-- d1832d
	sted1832d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1832d,
			Enable=>Enabled1832d,
			match=>matchd1832d,
			run=>run);

	Enabled1832d <= matchd1831d;
	-- d1833d
	sted1833d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1833d,
			Enable=>Enabled1833d,
			match=>matchd1833d,
			run=>run);

	-- d1834d
	sted1834d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1834d,
			Enable=>Enabled1834d,
			match=>matchd1834d,
			run=>run);

	Enabled1834d <= matchd1833d OR matchd1834d;
	-- d1835d
	sted1835d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1835d,
			Enable=>Enabled1835d,
			match=>matchd1835d,
			run=>run);

	Enabled1835d <= matchd1834d;
	-- d1836d
	sted1836d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1836d,
			Enable=>Enabled1836d,
			match=>matchd1836d,
			run=>run);

	Enabled1836d <= matchd1835d;
	-- d1837d
	sted1837d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1837d,
			Enable=>Enabled1837d,
			match=>matchd1837d,
			run=>run);

	Enabled1837d <= matchd1836d;
	-- d1838d
	sted1838d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1838d,
			Enable=>Enabled1838d,
			match=>matchd1838d,
			run=>run);

	Enabled1838d <= matchd1837d;
	-- d1839d
	sted1839d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1839d,
			Enable=>Enabled1839d,
			match=>matchd1839d,
			run=>run);

	Enabled1839d <= matchd1838d OR matchd1839d;
	-- d1840d
	sted1840d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1840d,
			Enable=>Enabled1840d,
			match=>matchd1840d,
			run=>run);

	Enabled1840d <= matchd1839d;
	-- d1841d
	sted1841d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1841d,
			Enable=>Enabled1841d,
			match=>matchd1841d,
			run=>run);

	Enabled1841d <= matchd1841d OR matchd1840d;
	-- d1842d
	sted1842d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1842d,
			Enable=>Enabled1842d,
			match=>matchd1842d,
			run=>run);

	Enabled1842d <= matchd1841d;
	-- d1843d
	sted1843d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1843d,
			Enable=>Enabled1843d,
			match=>matchd1843d,
			run=>run);

	Enabled1843d <= matchd1842d OR matchd1843d;
	-- d1844d
	sted1844d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1844d,
			Enable=>Enabled1844d,
			match=>matchd1844d,
			run=>run);

	Enabled1844d <= matchd1843d;
	-- d1845d
	sted1845d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1845d,
			Enable=>Enabled1845d,
			match=>matchd1845d,
			run=>run);

	Enabled1845d <= matchd1844d OR matchd1845d;
	-- d1846d
	sted1846d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1846d,
			Enable=>Enabled1846d,
			match=>matchd1846d,
			run=>run);

	Enabled1846d <= matchd1845d;
	-- d1847d
	sted1847d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1847d,
			Enable=>Enabled1847d,
			match=>matchd1847d,
			run=>run);

	Enabled1847d <= matchd1847d OR matchd1846d;
	-- d1848d
	sted1848d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1848d,
			Enable=>Enabled1848d,
			match=>matchd1848d,
			run=>run);

	Enabled1848d <= matchd1847d;
	-- d1849d
	sted1849d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1849d,
			Enable=>Enabled1849d,
			match=>matchd1849d,
			run=>run);

	Enabled1849d <= matchd1848d;
	-- d1850d
	sted1850d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1850d,
			Enable=>Enabled1850d,
			match=>matchd1850d,
			run=>run);

	Enabled1850d <= matchd1849d;
	-- d1852d
	sted1852d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1852d,
			Enable=>Enabled1852d,
			match=>matchd1852d,
			run=>run);

	-- d1853d
	sted1853d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1853d,
			Enable=>Enabled1853d,
			match=>matchd1853d,
			run=>run);

	Enabled1853d <= matchd1853d OR matchd1852d;
	-- d1854d
	sted1854d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1854d,
			Enable=>Enabled1854d,
			match=>matchd1854d,
			run=>run);

	Enabled1854d <= matchd1853d;
	-- d1855d
	sted1855d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1855d,
			Enable=>Enabled1855d,
			match=>matchd1855d,
			run=>run);

	Enabled1855d <= matchd1854d;
	-- d1856d
	sted1856d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1856d,
			Enable=>Enabled1856d,
			match=>matchd1856d,
			run=>run);

	Enabled1856d <= matchd1855d;
	-- d1857d
	sted1857d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1857d,
			Enable=>Enabled1857d,
			match=>matchd1857d,
			run=>run);

	Enabled1857d <= matchd1856d;
	-- d1858d
	sted1858d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1858d,
			Enable=>Enabled1858d,
			match=>matchd1858d,
			run=>run);

	Enabled1858d <= matchd1858d OR matchd1857d;
	-- d1859d
	sted1859d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1859d,
			Enable=>Enabled1859d,
			match=>matchd1859d,
			run=>run);

	Enabled1859d <= matchd1858d;
	-- d1860d
	sted1860d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1860d,
			Enable=>Enabled1860d,
			match=>matchd1860d,
			run=>run);

	Enabled1860d <= matchd1859d;
	-- d1861d
	sted1861d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1861d,
			Enable=>Enabled1861d,
			match=>matchd1861d,
			run=>run);

	Enabled1861d <= matchd1860d;
	-- d1862d
	sted1862d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1862d,
			Enable=>Enabled1862d,
			match=>matchd1862d,
			run=>run);

	reports(91) <= matchd1862d;
	Enabled1862d <= matchd1861d;
	-- d1863d
	sted1863d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1863d,
			Enable=>Enabled1863d,
			match=>matchd1863d,
			run=>run);

	-- d1864d
	sted1864d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1864d,
			Enable=>Enabled1864d,
			match=>matchd1864d,
			run=>run);

	Enabled1864d <= matchd1864d OR matchd1863d;
	-- d1865d
	sted1865d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1865d,
			Enable=>Enabled1865d,
			match=>matchd1865d,
			run=>run);

	Enabled1865d <= matchd1864d;
	-- d1866d
	sted1866d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1866d,
			Enable=>Enabled1866d,
			match=>matchd1866d,
			run=>run);

	Enabled1866d <= matchd1865d;
	-- d1867d
	sted1867d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1867d,
			Enable=>Enabled1867d,
			match=>matchd1867d,
			run=>run);

	Enabled1867d <= matchd1866d;
	-- d1868d
	sted1868d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1868d,
			Enable=>Enabled1868d,
			match=>matchd1868d,
			run=>run);

	Enabled1868d <= matchd1867d;
	-- d1869d
	sted1869d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1869d,
			Enable=>Enabled1869d,
			match=>matchd1869d,
			run=>run);

	Enabled1869d <= matchd1869d OR matchd1868d;
	-- d1870d
	sted1870d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1870d,
			Enable=>Enabled1870d,
			match=>matchd1870d,
			run=>run);

	Enabled1870d <= matchd1869d;
	-- d1871d
	sted1871d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1871d,
			Enable=>Enabled1871d,
			match=>matchd1871d,
			run=>run);

	Enabled1871d <= matchd1870d;
	-- d1872d
	sted1872d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1872d,
			Enable=>Enabled1872d,
			match=>matchd1872d,
			run=>run);

	Enabled1872d <= matchd1871d;
	-- d1873d
	sted1873d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1873d,
			Enable=>Enabled1873d,
			match=>matchd1873d,
			run=>run);

	Enabled1873d <= matchd1872d;
	-- d1874d
	sted1874d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1874d,
			Enable=>Enabled1874d,
			match=>matchd1874d,
			run=>run);

	reports(92) <= matchd1874d;
	Enabled1874d <= matchd1873d;
	-- d1875d
	sted1875d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1875d,
			Enable=>Enabled1875d,
			match=>matchd1875d,
			run=>run);

	-- d1876d
	sted1876d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1876d,
			Enable=>Enabled1876d,
			match=>matchd1876d,
			run=>run);

	Enabled1876d <= matchd1875d;
	-- d1877d
	sted1877d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1877d,
			Enable=>Enabled1877d,
			match=>matchd1877d,
			run=>run);

	Enabled1877d <= matchd1876d;
	-- d1878d
	sted1878d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1878d,
			Enable=>Enabled1878d,
			match=>matchd1878d,
			run=>run);

	Enabled1878d <= matchd1877d;
	-- d1879d
	sted1879d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1879d,
			Enable=>Enabled1879d,
			match=>matchd1879d,
			run=>run);

	Enabled1879d <= matchd1878d;
	-- d1880d
	sted1880d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1880d,
			Enable=>Enabled1880d,
			match=>matchd1880d,
			run=>run);

	Enabled1880d <= matchd1879d;
	-- d1881d
	sted1881d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1881d,
			Enable=>Enabled1881d,
			match=>matchd1881d,
			run=>run);

	Enabled1881d <= matchd1880d;
	-- d1882d
	sted1882d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1882d,
			Enable=>Enabled1882d,
			match=>matchd1882d,
			run=>run);

	Enabled1882d <= matchd1881d;
	-- d1883d
	sted1883d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1883d,
			Enable=>Enabled1883d,
			match=>matchd1883d,
			run=>run);

	Enabled1883d <= matchd1882d;
	-- d1884d
	sted1884d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1884d,
			Enable=>Enabled1884d,
			match=>matchd1884d,
			run=>run);

	Enabled1884d <= matchd1883d OR matchd1884d;
	-- d1885d
	sted1885d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1885d,
			Enable=>Enabled1885d,
			match=>matchd1885d,
			run=>run);

	Enabled1885d <= matchd1884d;
	-- d1886d
	sted1886d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1886d,
			Enable=>Enabled1886d,
			match=>matchd1886d,
			run=>run);

	Enabled1886d <= matchd1885d;
	-- d1887d
	sted1887d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1887d,
			Enable=>Enabled1887d,
			match=>matchd1887d,
			run=>run);

	Enabled1887d <= matchd1886d;
	-- d1888d
	sted1888d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1888d,
			Enable=>Enabled1888d,
			match=>matchd1888d,
			run=>run);

	reports(93) <= matchd1888d;
	Enabled1888d <= matchd1887d;
	-- d1889d
	sted1889d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1889d,
			Enable=>Enabled1889d,
			match=>matchd1889d,
			run=>run);

	-- d1890d
	sted1890d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1890d,
			Enable=>Enabled1890d,
			match=>matchd1890d,
			run=>run);

	Enabled1890d <= matchd1890d OR matchd1889d;
	-- d1891d
	sted1891d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1891d,
			Enable=>Enabled1891d,
			match=>matchd1891d,
			run=>run);

	Enabled1891d <= matchd1890d;
	-- d1892d
	sted1892d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1892d,
			Enable=>Enabled1892d,
			match=>matchd1892d,
			run=>run);

	Enabled1892d <= matchd1891d;
	-- d1893d
	sted1893d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1893d,
			Enable=>Enabled1893d,
			match=>matchd1893d,
			run=>run);

	Enabled1893d <= matchd1892d;
	-- d1894d
	sted1894d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1894d,
			Enable=>Enabled1894d,
			match=>matchd1894d,
			run=>run);

	Enabled1894d <= matchd1893d;
	-- d1895d
	sted1895d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1895d,
			Enable=>Enabled1895d,
			match=>matchd1895d,
			run=>run);

	Enabled1895d <= matchd1894d OR matchd1895d;
	-- d1896d
	sted1896d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1896d,
			Enable=>Enabled1896d,
			match=>matchd1896d,
			run=>run);

	Enabled1896d <= matchd1895d;
	-- d1897d
	sted1897d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1897d,
			Enable=>Enabled1897d,
			match=>matchd1897d,
			run=>run);

	Enabled1897d <= matchd1896d;
	-- d1898d
	sted1898d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1898d,
			Enable=>Enabled1898d,
			match=>matchd1898d,
			run=>run);

	Enabled1898d <= matchd1897d;
	-- d1899d
	sted1899d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1899d,
			Enable=>Enabled1899d,
			match=>matchd1899d,
			run=>run);

	Enabled1899d <= matchd1898d;
	-- d1900d
	sted1900d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1900d,
			Enable=>Enabled1900d,
			match=>matchd1900d,
			run=>run);

	Enabled1900d <= matchd1900d OR matchd1899d;
	-- d1901d
	sted1901d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1901d,
			Enable=>Enabled1901d,
			match=>matchd1901d,
			run=>run);

	Enabled1901d <= matchd1900d;
	-- d1902d
	sted1902d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1902d,
			Enable=>Enabled1902d,
			match=>matchd1902d,
			run=>run);

	Enabled1902d <= matchd1901d;
	-- d1903d
	sted1903d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1903d,
			Enable=>Enabled1903d,
			match=>matchd1903d,
			run=>run);

	Enabled1903d <= matchd1902d;
	-- d1904d
	sted1904d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1904d,
			Enable=>Enabled1904d,
			match=>matchd1904d,
			run=>run);

	reports(94) <= matchd1904d;
	Enabled1904d <= matchd1903d;
	-- d1905d
	sted1905d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1905d,
			Enable=>Enabled1905d,
			match=>matchd1905d,
			run=>run);

	-- d1906d
	sted1906d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1906d,
			Enable=>Enabled1906d,
			match=>matchd1906d,
			run=>run);

	Enabled1906d <= matchd1905d OR matchd1906d;
	-- d1907d
	sted1907d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1907d,
			Enable=>Enabled1907d,
			match=>matchd1907d,
			run=>run);

	Enabled1907d <= matchd1906d;
	-- d1908d
	sted1908d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1908d,
			Enable=>Enabled1908d,
			match=>matchd1908d,
			run=>run);

	Enabled1908d <= matchd1907d;
	-- d1909d
	sted1909d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1909d,
			Enable=>Enabled1909d,
			match=>matchd1909d,
			run=>run);

	Enabled1909d <= matchd1908d;
	-- d1910d
	sted1910d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1910d,
			Enable=>Enabled1910d,
			match=>matchd1910d,
			run=>run);

	Enabled1910d <= matchd1909d;
	-- d1911d
	sted1911d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1911d,
			Enable=>Enabled1911d,
			match=>matchd1911d,
			run=>run);

	Enabled1911d <= matchd1911d OR matchd1910d;
	-- d1912d
	sted1912d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1912d,
			Enable=>Enabled1912d,
			match=>matchd1912d,
			run=>run);

	Enabled1912d <= matchd1911d;
	-- d1913d
	sted1913d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1913d,
			Enable=>Enabled1913d,
			match=>matchd1913d,
			run=>run);

	Enabled1913d <= matchd1912d;
	-- d1914d
	sted1914d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1914d,
			Enable=>Enabled1914d,
			match=>matchd1914d,
			run=>run);

	Enabled1914d <= matchd1913d;
	-- d1915d
	sted1915d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1915d,
			Enable=>Enabled1915d,
			match=>matchd1915d,
			run=>run);

	Enabled1915d <= matchd1914d;
	-- d1916d
	sted1916d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1916d,
			Enable=>Enabled1916d,
			match=>matchd1916d,
			run=>run);

	reports(95) <= matchd1916d;
	Enabled1916d <= matchd1915d;
	-- d1917d
	sted1917d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1917d,
			Enable=>Enabled1917d,
			match=>matchd1917d,
			run=>run);

	-- d1918d
	sted1918d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1918d,
			Enable=>Enabled1918d,
			match=>matchd1918d,
			run=>run);

	Enabled1918d <= matchd1917d OR matchd1918d;
	-- d1919d
	sted1919d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1919d,
			Enable=>Enabled1919d,
			match=>matchd1919d,
			run=>run);

	Enabled1919d <= matchd1918d;
	-- d1920d
	sted1920d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1920d,
			Enable=>Enabled1920d,
			match=>matchd1920d,
			run=>run);

	Enabled1920d <= matchd1919d;
	-- d1921d
	sted1921d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1921d,
			Enable=>Enabled1921d,
			match=>matchd1921d,
			run=>run);

	Enabled1921d <= matchd1920d;
	-- d1922d
	sted1922d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1922d,
			Enable=>Enabled1922d,
			match=>matchd1922d,
			run=>run);

	Enabled1922d <= matchd1921d;
	-- d1923d
	sted1923d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1923d,
			Enable=>Enabled1923d,
			match=>matchd1923d,
			run=>run);

	Enabled1923d <= matchd1922d;
	-- d1924d
	sted1924d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1924d,
			Enable=>Enabled1924d,
			match=>matchd1924d,
			run=>run);

	Enabled1924d <= matchd1923d OR matchd1924d;
	-- d1925d
	sted1925d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1925d,
			Enable=>Enabled1925d,
			match=>matchd1925d,
			run=>run);

	Enabled1925d <= matchd1924d;
	-- d1926d
	sted1926d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1926d,
			Enable=>Enabled1926d,
			match=>matchd1926d,
			run=>run);

	Enabled1926d <= matchd1925d;
	-- d1927d
	sted1927d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1927d,
			Enable=>Enabled1927d,
			match=>matchd1927d,
			run=>run);

	Enabled1927d <= matchd1926d;
	-- d1928d
	sted1928d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1928d,
			Enable=>Enabled1928d,
			match=>matchd1928d,
			run=>run);

	Enabled1928d <= matchd1927d;
	-- d1929d
	sted1929d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1929d,
			Enable=>Enabled1929d,
			match=>matchd1929d,
			run=>run);

	Enabled1929d <= matchd1928d;
	-- d1930d
	sted1930d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1930d,
			Enable=>Enabled1930d,
			match=>matchd1930d,
			run=>run);

	Enabled1930d <= matchd1930d OR matchd1929d;
	-- d1931d
	sted1931d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1931d,
			Enable=>Enabled1931d,
			match=>matchd1931d,
			run=>run);

	Enabled1931d <= matchd1930d;
	-- d1932d
	sted1932d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1932d,
			Enable=>Enabled1932d,
			match=>matchd1932d,
			run=>run);

	Enabled1932d <= matchd1931d;
	-- d1933d
	sted1933d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1933d,
			Enable=>Enabled1933d,
			match=>matchd1933d,
			run=>run);

	Enabled1933d <= matchd1932d;
	-- d1934d
	sted1934d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1934d,
			Enable=>Enabled1934d,
			match=>matchd1934d,
			run=>run);

	reports(96) <= matchd1934d;
	Enabled1934d <= matchd1933d;
	-- d1935d
	sted1935d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1935d,
			Enable=>Enabled1935d,
			match=>matchd1935d,
			run=>run);

	-- d1936d
	sted1936d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1936d,
			Enable=>Enabled1936d,
			match=>matchd1936d,
			run=>run);

	Enabled1936d <= matchd1936d OR matchd1935d;
	-- d1937d
	sted1937d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1937d,
			Enable=>Enabled1937d,
			match=>matchd1937d,
			run=>run);

	Enabled1937d <= matchd1936d;
	-- d1938d
	sted1938d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1938d,
			Enable=>Enabled1938d,
			match=>matchd1938d,
			run=>run);

	Enabled1938d <= matchd1937d;
	-- d1939d
	sted1939d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1939d,
			Enable=>Enabled1939d,
			match=>matchd1939d,
			run=>run);

	Enabled1939d <= matchd1938d;
	-- d1940d
	sted1940d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1940d,
			Enable=>Enabled1940d,
			match=>matchd1940d,
			run=>run);

	Enabled1940d <= matchd1939d;
	-- d1941d
	sted1941d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1941d,
			Enable=>Enabled1941d,
			match=>matchd1941d,
			run=>run);

	Enabled1941d <= matchd1940d OR matchd1941d;
	-- d1942d
	sted1942d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1942d,
			Enable=>Enabled1942d,
			match=>matchd1942d,
			run=>run);

	Enabled1942d <= matchd1941d;
	-- d1943d
	sted1943d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1943d,
			Enable=>Enabled1943d,
			match=>matchd1943d,
			run=>run);

	Enabled1943d <= matchd1942d;
	-- d1944d
	sted1944d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1944d,
			Enable=>Enabled1944d,
			match=>matchd1944d,
			run=>run);

	reports(97) <= matchd1944d;
	Enabled1944d <= matchd1943d;
	-- d1945d
	sted1945d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1945d,
			Enable=>Enabled1945d,
			match=>matchd1945d,
			run=>run);

	-- d1946d
	sted1946d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1946d,
			Enable=>Enabled1946d,
			match=>matchd1946d,
			run=>run);

	Enabled1946d <= matchd1946d OR matchd1945d;
	-- d1947d
	sted1947d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1947d,
			Enable=>Enabled1947d,
			match=>matchd1947d,
			run=>run);

	Enabled1947d <= matchd1946d;
	-- d1948d
	sted1948d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1948d,
			Enable=>Enabled1948d,
			match=>matchd1948d,
			run=>run);

	Enabled1948d <= matchd1947d;
	-- d1949d
	sted1949d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1949d,
			Enable=>Enabled1949d,
			match=>matchd1949d,
			run=>run);

	Enabled1949d <= matchd1948d;
	-- d1950d
	sted1950d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1950d,
			Enable=>Enabled1950d,
			match=>matchd1950d,
			run=>run);

	Enabled1950d <= matchd1949d;
	-- d1951d
	sted1951d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1951d,
			Enable=>Enabled1951d,
			match=>matchd1951d,
			run=>run);

	Enabled1951d <= matchd1950d;
	-- d1952d
	sted1952d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1952d,
			Enable=>Enabled1952d,
			match=>matchd1952d,
			run=>run);

	Enabled1952d <= matchd1951d OR matchd1952d;
	-- d1953d
	sted1953d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1953d,
			Enable=>Enabled1953d,
			match=>matchd1953d,
			run=>run);

	Enabled1953d <= matchd1952d;
	-- d1954d
	sted1954d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1954d,
			Enable=>Enabled1954d,
			match=>matchd1954d,
			run=>run);

	Enabled1954d <= matchd1953d;
	-- d1955d
	sted1955d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1955d,
			Enable=>Enabled1955d,
			match=>matchd1955d,
			run=>run);

	Enabled1955d <= matchd1954d;
	-- d1956d
	sted1956d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1956d,
			Enable=>Enabled1956d,
			match=>matchd1956d,
			run=>run);

	reports(98) <= matchd1956d;
	Enabled1956d <= matchd1955d;
	-- d1957d
	sted1957d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1957d,
			Enable=>Enabled1957d,
			match=>matchd1957d,
			run=>run);

	-- d1958d
	sted1958d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1958d,
			Enable=>Enabled1958d,
			match=>matchd1958d,
			run=>run);

	Enabled1958d <= matchd1957d OR matchd1958d;
	-- d1959d
	sted1959d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1959d,
			Enable=>Enabled1959d,
			match=>matchd1959d,
			run=>run);

	Enabled1959d <= matchd1958d;
	-- d1960d
	sted1960d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1960d,
			Enable=>Enabled1960d,
			match=>matchd1960d,
			run=>run);

	Enabled1960d <= matchd1959d;
	-- d1961d
	sted1961d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1961d,
			Enable=>Enabled1961d,
			match=>matchd1961d,
			run=>run);

	Enabled1961d <= matchd1960d;
	-- d1962d
	sted1962d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1962d,
			Enable=>Enabled1962d,
			match=>matchd1962d,
			run=>run);

	Enabled1962d <= matchd1961d;
	-- d1963d
	sted1963d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1963d,
			Enable=>Enabled1963d,
			match=>matchd1963d,
			run=>run);

	Enabled1963d <= matchd1962d OR matchd1963d;
	-- d1964d
	sted1964d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1964d,
			Enable=>Enabled1964d,
			match=>matchd1964d,
			run=>run);

	Enabled1964d <= matchd1963d;
	-- d1965d
	sted1965d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1965d,
			Enable=>Enabled1965d,
			match=>matchd1965d,
			run=>run);

	Enabled1965d <= matchd1964d;
	-- d1966d
	sted1966d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1966d,
			Enable=>Enabled1966d,
			match=>matchd1966d,
			run=>run);

	Enabled1966d <= matchd1965d;
	-- d1967d
	sted1967d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1967d,
			Enable=>Enabled1967d,
			match=>matchd1967d,
			run=>run);

	Enabled1967d <= matchd1966d;
	-- d1968d
	sted1968d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1968d,
			Enable=>Enabled1968d,
			match=>matchd1968d,
			run=>run);

	reports(99) <= matchd1968d;
	Enabled1968d <= matchd1967d;
	-- d1969d
	sted1969d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1969d,
			Enable=>Enabled1969d,
			match=>matchd1969d,
			run=>run);

	-- d1970d
	sted1970d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1970d,
			Enable=>Enabled1970d,
			match=>matchd1970d,
			run=>run);

	Enabled1970d <= matchd1969d OR matchd1970d;
	-- d1971d
	sted1971d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1971d,
			Enable=>Enabled1971d,
			match=>matchd1971d,
			run=>run);

	Enabled1971d <= matchd1970d;
	-- d1972d
	sted1972d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1972d,
			Enable=>Enabled1972d,
			match=>matchd1972d,
			run=>run);

	Enabled1972d <= matchd1971d;
	-- d1973d
	sted1973d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1973d,
			Enable=>Enabled1973d,
			match=>matchd1973d,
			run=>run);

	Enabled1973d <= matchd1972d;
	-- d1974d
	sted1974d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1974d,
			Enable=>Enabled1974d,
			match=>matchd1974d,
			run=>run);

	Enabled1974d <= matchd1973d;
	-- d1975d
	sted1975d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1975d,
			Enable=>Enabled1975d,
			match=>matchd1975d,
			run=>run);

	Enabled1975d <= matchd1975d OR matchd1974d;
	-- d1976d
	sted1976d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1976d,
			Enable=>Enabled1976d,
			match=>matchd1976d,
			run=>run);

	Enabled1976d <= matchd1975d;
	-- d1977d
	sted1977d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1977d,
			Enable=>Enabled1977d,
			match=>matchd1977d,
			run=>run);

	Enabled1977d <= matchd1976d;
	-- d1978d
	sted1978d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1978d,
			Enable=>Enabled1978d,
			match=>matchd1978d,
			run=>run);

	Enabled1978d <= matchd1977d;
	-- d1979d
	sted1979d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1979d,
			Enable=>Enabled1979d,
			match=>matchd1979d,
			run=>run);

	Enabled1979d <= matchd1978d;
	-- d1980d
	sted1980d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1980d,
			Enable=>Enabled1980d,
			match=>matchd1980d,
			run=>run);

	reports(100) <= matchd1980d;
	Enabled1980d <= matchd1979d;
	-- d1981d
	sted1981d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1981d,
			Enable=>Enabled1981d,
			match=>matchd1981d,
			run=>run);

	-- d1982d
	sted1982d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1982d,
			Enable=>Enabled1982d,
			match=>matchd1982d,
			run=>run);

	Enabled1982d <= matchd1982d OR matchd1981d;
	-- d1983d
	sted1983d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1983d,
			Enable=>Enabled1983d,
			match=>matchd1983d,
			run=>run);

	Enabled1983d <= matchd1982d;
	-- d1984d
	sted1984d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1984d,
			Enable=>Enabled1984d,
			match=>matchd1984d,
			run=>run);

	Enabled1984d <= matchd1983d;
	-- d1985d
	sted1985d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1985d,
			Enable=>Enabled1985d,
			match=>matchd1985d,
			run=>run);

	Enabled1985d <= matchd1984d;
	-- d1986d
	sted1986d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1986d,
			Enable=>Enabled1986d,
			match=>matchd1986d,
			run=>run);

	Enabled1986d <= matchd1985d;
	-- d1987d
	sted1987d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1987d,
			Enable=>Enabled1987d,
			match=>matchd1987d,
			run=>run);

	Enabled1987d <= matchd1986d OR matchd1987d;
	-- d1988d
	sted1988d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1988d,
			Enable=>Enabled1988d,
			match=>matchd1988d,
			run=>run);

	Enabled1988d <= matchd1987d;
	-- d1989d
	sted1989d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1989d,
			Enable=>Enabled1989d,
			match=>matchd1989d,
			run=>run);

	Enabled1989d <= matchd1988d;
	-- d1990d
	sted1990d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1990d,
			Enable=>Enabled1990d,
			match=>matchd1990d,
			run=>run);

	Enabled1990d <= matchd1989d;
	-- d1991d
	sted1991d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1991d,
			Enable=>Enabled1991d,
			match=>matchd1991d,
			run=>run);

	Enabled1991d <= matchd1990d;
	-- d1992d
	sted1992d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1992d,
			Enable=>Enabled1992d,
			match=>matchd1992d,
			run=>run);

	Enabled1992d <= matchd1991d OR matchd1992d;
	-- d1993d
	sted1993d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1993d,
			Enable=>Enabled1993d,
			match=>matchd1993d,
			run=>run);

	Enabled1993d <= matchd1992d;
	-- d1994d
	sted1994d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1994d,
			Enable=>Enabled1994d,
			match=>matchd1994d,
			run=>run);

	Enabled1994d <= matchd1993d;
	-- d1995d
	sted1995d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1995d,
			Enable=>Enabled1995d,
			match=>matchd1995d,
			run=>run);

	reports(101) <= matchd1995d;
	Enabled1995d <= matchd1994d;
	-- d1996d
	sted1996d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1996d,
			Enable=>Enabled1996d,
			match=>matchd1996d,
			run=>run);

	-- d1997d
	sted1997d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1997d,
			Enable=>Enabled1997d,
			match=>matchd1997d,
			run=>run);

	Enabled1997d <= matchd1997d OR matchd1996d;
	-- d1998d
	sted1998d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1998d,
			Enable=>Enabled1998d,
			match=>matchd1998d,
			run=>run);

	Enabled1998d <= matchd1997d;
	-- d1999d
	sted1999d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord1999d,
			Enable=>Enabled1999d,
			match=>matchd1999d,
			run=>run);

	Enabled1999d <= matchd1998d;
	-- d2000d
	sted2000d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2000d,
			Enable=>Enabled2000d,
			match=>matchd2000d,
			run=>run);

	Enabled2000d <= matchd1999d;
	-- d2001d
	sted2001d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2001d,
			Enable=>Enabled2001d,
			match=>matchd2001d,
			run=>run);

	Enabled2001d <= matchd2000d;
	-- d2002d
	sted2002d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2002d,
			Enable=>Enabled2002d,
			match=>matchd2002d,
			run=>run);

	Enabled2002d <= matchd2001d;
	-- d2003d
	sted2003d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2003d,
			Enable=>Enabled2003d,
			match=>matchd2003d,
			run=>run);

	Enabled2003d <= matchd2002d OR matchd2003d;
	-- d2004d
	sted2004d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2004d,
			Enable=>Enabled2004d,
			match=>matchd2004d,
			run=>run);

	Enabled2004d <= matchd2003d;
	-- d2005d
	sted2005d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2005d,
			Enable=>Enabled2005d,
			match=>matchd2005d,
			run=>run);

	Enabled2005d <= matchd2004d;
	-- d2006d
	sted2006d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2006d,
			Enable=>Enabled2006d,
			match=>matchd2006d,
			run=>run);

	Enabled2006d <= matchd2005d;
	-- d2007d
	sted2007d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2007d,
			Enable=>Enabled2007d,
			match=>matchd2007d,
			run=>run);

	Enabled2007d <= matchd2006d;
	-- d2008d
	sted2008d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2008d,
			Enable=>Enabled2008d,
			match=>matchd2008d,
			run=>run);

	Enabled2008d <= matchd2007d OR matchd2008d;
	-- d2009d
	sted2009d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2009d,
			Enable=>Enabled2009d,
			match=>matchd2009d,
			run=>run);

	Enabled2009d <= matchd2008d;
	-- d2010d
	sted2010d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2010d,
			Enable=>Enabled2010d,
			match=>matchd2010d,
			run=>run);

	Enabled2010d <= matchd2009d;
	-- d2011d
	sted2011d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2011d,
			Enable=>Enabled2011d,
			match=>matchd2011d,
			run=>run);

	Enabled2011d <= matchd2010d;
	-- d2012d
	sted2012d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2012d,
			Enable=>Enabled2012d,
			match=>matchd2012d,
			run=>run);

	Enabled2012d <= matchd2011d;
	-- d2013d
	sted2013d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2013d,
			Enable=>Enabled2013d,
			match=>matchd2013d,
			run=>run);

	reports(102) <= matchd2013d;
	Enabled2013d <= matchd2012d;
	-- d2014d
	sted2014d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2014d,
			Enable=>Enabled2014d,
			match=>matchd2014d,
			run=>run);

	-- d2015d
	sted2015d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2015d,
			Enable=>Enabled2015d,
			match=>matchd2015d,
			run=>run);

	Enabled2015d <= matchd2015d OR matchd2014d;
	-- d2016d
	sted2016d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2016d,
			Enable=>Enabled2016d,
			match=>matchd2016d,
			run=>run);

	Enabled2016d <= matchd2015d;
	-- d2017d
	sted2017d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2017d,
			Enable=>Enabled2017d,
			match=>matchd2017d,
			run=>run);

	Enabled2017d <= matchd2016d;
	-- d2018d
	sted2018d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2018d,
			Enable=>Enabled2018d,
			match=>matchd2018d,
			run=>run);

	Enabled2018d <= matchd2017d;
	-- d2019d
	sted2019d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2019d,
			Enable=>Enabled2019d,
			match=>matchd2019d,
			run=>run);

	Enabled2019d <= matchd2018d;
	-- d2020d
	sted2020d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2020d,
			Enable=>Enabled2020d,
			match=>matchd2020d,
			run=>run);

	Enabled2020d <= matchd2020d OR matchd2019d;
	-- d2021d
	sted2021d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2021d,
			Enable=>Enabled2021d,
			match=>matchd2021d,
			run=>run);

	Enabled2021d <= matchd2020d;
	-- d2022d
	sted2022d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2022d,
			Enable=>Enabled2022d,
			match=>matchd2022d,
			run=>run);

	Enabled2022d <= matchd2021d;
	-- d2023d
	sted2023d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2023d,
			Enable=>Enabled2023d,
			match=>matchd2023d,
			run=>run);

	Enabled2023d <= matchd2022d;
	-- d2024d
	sted2024d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2024d,
			Enable=>Enabled2024d,
			match=>matchd2024d,
			run=>run);

	Enabled2024d <= matchd2023d;
	-- d2025d
	sted2025d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2025d,
			Enable=>Enabled2025d,
			match=>matchd2025d,
			run=>run);

	reports(103) <= matchd2025d;
	Enabled2025d <= matchd2024d;
	-- d2026d
	sted2026d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2026d,
			Enable=>Enabled2026d,
			match=>matchd2026d,
			run=>run);

	-- d2027d
	sted2027d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2027d,
			Enable=>Enabled2027d,
			match=>matchd2027d,
			run=>run);

	Enabled2027d <= matchd2026d;
	-- d2028d
	sted2028d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2028d,
			Enable=>Enabled2028d,
			match=>matchd2028d,
			run=>run);

	Enabled2028d <= matchd2027d;
	-- d2029d
	sted2029d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2029d,
			Enable=>Enabled2029d,
			match=>matchd2029d,
			run=>run);

	Enabled2029d <= matchd2028d;
	-- d2030d
	sted2030d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2030d,
			Enable=>Enabled2030d,
			match=>matchd2030d,
			run=>run);

	Enabled2030d <= matchd2029d;
	-- d2031d
	sted2031d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2031d,
			Enable=>Enabled2031d,
			match=>matchd2031d,
			run=>run);

	Enabled2031d <= matchd2030d;
	-- d2032d
	sted2032d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2032d,
			Enable=>Enabled2032d,
			match=>matchd2032d,
			run=>run);

	Enabled2032d <= matchd2031d;
	-- d2033d
	sted2033d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2033d,
			Enable=>Enabled2033d,
			match=>matchd2033d,
			run=>run);

	Enabled2033d <= matchd2032d OR matchd2033d;
	-- d2034d
	sted2034d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2034d,
			Enable=>Enabled2034d,
			match=>matchd2034d,
			run=>run);

	Enabled2034d <= matchd2033d;
	-- d2035d
	sted2035d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2035d,
			Enable=>Enabled2035d,
			match=>matchd2035d,
			run=>run);

	Enabled2035d <= matchd2034d;
	-- d2036d
	sted2036d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2036d,
			Enable=>Enabled2036d,
			match=>matchd2036d,
			run=>run);

	Enabled2036d <= matchd2035d;
	-- d2037d
	sted2037d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2037d,
			Enable=>Enabled2037d,
			match=>matchd2037d,
			run=>run);

	reports(104) <= matchd2037d;
	Enabled2037d <= matchd2036d;
	-- d2038d
	sted2038d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2038d,
			Enable=>Enabled2038d,
			match=>matchd2038d,
			run=>run);

	-- d2039d
	sted2039d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2039d,
			Enable=>Enabled2039d,
			match=>matchd2039d,
			run=>run);

	Enabled2039d <= matchd2039d OR matchd2038d;
	-- d2040d
	sted2040d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2040d,
			Enable=>Enabled2040d,
			match=>matchd2040d,
			run=>run);

	Enabled2040d <= matchd2039d;
	-- d2041d
	sted2041d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2041d,
			Enable=>Enabled2041d,
			match=>matchd2041d,
			run=>run);

	Enabled2041d <= matchd2040d;
	-- d2042d
	sted2042d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2042d,
			Enable=>Enabled2042d,
			match=>matchd2042d,
			run=>run);

	Enabled2042d <= matchd2041d;
	-- d2043d
	sted2043d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2043d,
			Enable=>Enabled2043d,
			match=>matchd2043d,
			run=>run);

	Enabled2043d <= matchd2042d;
	-- d2044d
	sted2044d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2044d,
			Enable=>Enabled2044d,
			match=>matchd2044d,
			run=>run);

	Enabled2044d <= matchd2044d OR matchd2043d;
	-- d2045d
	sted2045d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2045d,
			Enable=>Enabled2045d,
			match=>matchd2045d,
			run=>run);

	Enabled2045d <= matchd2044d;
	-- d2046d
	sted2046d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2046d,
			Enable=>Enabled2046d,
			match=>matchd2046d,
			run=>run);

	Enabled2046d <= matchd2045d;
	-- d2047d
	sted2047d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2047d,
			Enable=>Enabled2047d,
			match=>matchd2047d,
			run=>run);

	Enabled2047d <= matchd2046d;
	-- d2048d
	sted2048d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2048d,
			Enable=>Enabled2048d,
			match=>matchd2048d,
			run=>run);

	Enabled2048d <= matchd2047d;
	-- d2049d
	sted2049d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2049d,
			Enable=>Enabled2049d,
			match=>matchd2049d,
			run=>run);

	reports(105) <= matchd2049d;
	Enabled2049d <= matchd2048d;
	-- d2050d
	sted2050d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2050d,
			Enable=>Enabled2050d,
			match=>matchd2050d,
			run=>run);

	-- d2051d
	sted2051d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2051d,
			Enable=>Enabled2051d,
			match=>matchd2051d,
			run=>run);

	Enabled2051d <= matchd2050d;
	-- d2052d
	sted2052d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2052d,
			Enable=>Enabled2052d,
			match=>matchd2052d,
			run=>run);

	Enabled2052d <= matchd2051d;
	-- d2053d
	sted2053d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2053d,
			Enable=>Enabled2053d,
			match=>matchd2053d,
			run=>run);

	Enabled2053d <= matchd2052d;
	-- d2054d
	sted2054d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2054d,
			Enable=>Enabled2054d,
			match=>matchd2054d,
			run=>run);

	Enabled2054d <= matchd2053d;
	-- d2055d
	sted2055d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2055d,
			Enable=>Enabled2055d,
			match=>matchd2055d,
			run=>run);

	Enabled2055d <= matchd2054d;
	-- d2056d
	sted2056d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2056d,
			Enable=>Enabled2056d,
			match=>matchd2056d,
			run=>run);

	Enabled2056d <= matchd2055d;
	-- d2057d
	sted2057d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2057d,
			Enable=>Enabled2057d,
			match=>matchd2057d,
			run=>run);

	Enabled2057d <= matchd2056d;
	-- d2058d
	sted2058d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2058d,
			Enable=>Enabled2058d,
			match=>matchd2058d,
			run=>run);

	Enabled2058d <= matchd2057d;
	-- d2059d
	sted2059d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2059d,
			Enable=>Enabled2059d,
			match=>matchd2059d,
			run=>run);

	Enabled2059d <= matchd2058d;
	-- d2060d
	sted2060d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2060d,
			Enable=>Enabled2060d,
			match=>matchd2060d,
			run=>run);

	Enabled2060d <= matchd2060d OR matchd2059d;
	-- d2061d
	sted2061d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2061d,
			Enable=>Enabled2061d,
			match=>matchd2061d,
			run=>run);

	Enabled2061d <= matchd2060d;
	-- d2062d
	sted2062d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2062d,
			Enable=>Enabled2062d,
			match=>matchd2062d,
			run=>run);

	Enabled2062d <= matchd2061d;
	-- d2063d
	sted2063d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2063d,
			Enable=>Enabled2063d,
			match=>matchd2063d,
			run=>run);

	Enabled2063d <= matchd2062d;
	-- d2064d
	sted2064d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2064d,
			Enable=>Enabled2064d,
			match=>matchd2064d,
			run=>run);

	reports(106) <= matchd2064d;
	Enabled2064d <= matchd2063d;
	-- d2065d
	sted2065d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2065d,
			Enable=>Enabled2065d,
			match=>matchd2065d,
			run=>run);

	-- d2066d
	sted2066d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2066d,
			Enable=>Enabled2066d,
			match=>matchd2066d,
			run=>run);

	Enabled2066d <= matchd2065d;
	-- d2067d
	sted2067d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2067d,
			Enable=>Enabled2067d,
			match=>matchd2067d,
			run=>run);

	Enabled2067d <= matchd2066d;
	-- d2068d
	sted2068d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2068d,
			Enable=>Enabled2068d,
			match=>matchd2068d,
			run=>run);

	Enabled2068d <= matchd2067d;
	-- d2069d
	sted2069d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2069d,
			Enable=>Enabled2069d,
			match=>matchd2069d,
			run=>run);

	Enabled2069d <= matchd2068d;
	-- d2070d
	sted2070d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2070d,
			Enable=>Enabled2070d,
			match=>matchd2070d,
			run=>run);

	Enabled2070d <= matchd2069d;
	-- d2071d
	sted2071d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2071d,
			Enable=>Enabled2071d,
			match=>matchd2071d,
			run=>run);

	Enabled2071d <= matchd2070d;
	-- d2072d
	sted2072d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2072d,
			Enable=>Enabled2072d,
			match=>matchd2072d,
			run=>run);

	Enabled2072d <= matchd2071d;
	-- d2073d
	sted2073d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2073d,
			Enable=>Enabled2073d,
			match=>matchd2073d,
			run=>run);

	Enabled2073d <= matchd2072d;
	-- d2074d
	sted2074d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2074d,
			Enable=>Enabled2074d,
			match=>matchd2074d,
			run=>run);

	Enabled2074d <= matchd2073d;
	-- d2075d
	sted2075d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2075d,
			Enable=>Enabled2075d,
			match=>matchd2075d,
			run=>run);

	Enabled2075d <= matchd2075d OR matchd2074d;
	-- d2076d
	sted2076d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2076d,
			Enable=>Enabled2076d,
			match=>matchd2076d,
			run=>run);

	Enabled2076d <= matchd2075d;
	-- d2077d
	sted2077d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2077d,
			Enable=>Enabled2077d,
			match=>matchd2077d,
			run=>run);

	Enabled2077d <= matchd2076d;
	-- d2078d
	sted2078d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2078d,
			Enable=>Enabled2078d,
			match=>matchd2078d,
			run=>run);

	Enabled2078d <= matchd2077d;
	-- d2079d
	sted2079d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2079d,
			Enable=>Enabled2079d,
			match=>matchd2079d,
			run=>run);

	reports(107) <= matchd2079d;
	Enabled2079d <= matchd2078d;
	-- d2080d
	sted2080d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2080d,
			Enable=>Enabled2080d,
			match=>matchd2080d,
			run=>run);

	-- d2081d
	sted2081d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2081d,
			Enable=>Enabled2081d,
			match=>matchd2081d,
			run=>run);

	Enabled2081d <= matchd2080d OR matchd2081d;
	-- d2082d
	sted2082d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2082d,
			Enable=>Enabled2082d,
			match=>matchd2082d,
			run=>run);

	Enabled2082d <= matchd2081d;
	-- d2083d
	sted2083d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2083d,
			Enable=>Enabled2083d,
			match=>matchd2083d,
			run=>run);

	Enabled2083d <= matchd2082d;
	-- d2084d
	sted2084d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2084d,
			Enable=>Enabled2084d,
			match=>matchd2084d,
			run=>run);

	Enabled2084d <= matchd2083d;
	-- d2085d
	sted2085d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2085d,
			Enable=>Enabled2085d,
			match=>matchd2085d,
			run=>run);

	Enabled2085d <= matchd2084d;
	-- d2086d
	sted2086d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2086d,
			Enable=>Enabled2086d,
			match=>matchd2086d,
			run=>run);

	Enabled2086d <= matchd2085d;
	-- d2087d
	sted2087d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2087d,
			Enable=>Enabled2087d,
			match=>matchd2087d,
			run=>run);

	Enabled2087d <= matchd2086d;
	-- d2088d
	sted2088d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2088d,
			Enable=>Enabled2088d,
			match=>matchd2088d,
			run=>run);

	Enabled2088d <= matchd2087d;
	-- d2089d
	sted2089d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2089d,
			Enable=>Enabled2089d,
			match=>matchd2089d,
			run=>run);

	Enabled2089d <= matchd2088d;
	-- d2090d
	sted2090d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2090d,
			Enable=>Enabled2090d,
			match=>matchd2090d,
			run=>run);

	Enabled2090d <= matchd2089d;
	-- d2091d
	sted2091d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2091d,
			Enable=>Enabled2091d,
			match=>matchd2091d,
			run=>run);

	Enabled2091d <= matchd2090d;
	-- d2092d
	sted2092d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2092d,
			Enable=>Enabled2092d,
			match=>matchd2092d,
			run=>run);

	Enabled2092d <= matchd2091d;
	-- d2093d
	sted2093d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2093d,
			Enable=>Enabled2093d,
			match=>matchd2093d,
			run=>run);

	Enabled2093d <= matchd2092d;
	-- d2094d
	sted2094d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2094d,
			Enable=>Enabled2094d,
			match=>matchd2094d,
			run=>run);

	reports(108) <= matchd2094d;
	Enabled2094d <= matchd2093d;
	-- d2095d
	sted2095d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2095d,
			Enable=>Enabled2095d,
			match=>matchd2095d,
			run=>run);

	-- d2096d
	sted2096d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2096d,
			Enable=>Enabled2096d,
			match=>matchd2096d,
			run=>run);

	Enabled2096d <= matchd2095d OR matchd2096d;
	-- d2097d
	sted2097d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2097d,
			Enable=>Enabled2097d,
			match=>matchd2097d,
			run=>run);

	Enabled2097d <= matchd2096d;
	-- d2098d
	sted2098d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2098d,
			Enable=>Enabled2098d,
			match=>matchd2098d,
			run=>run);

	Enabled2098d <= matchd2097d;
	-- d2099d
	sted2099d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2099d,
			Enable=>Enabled2099d,
			match=>matchd2099d,
			run=>run);

	Enabled2099d <= matchd2098d;
	-- d2100d
	sted2100d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2100d,
			Enable=>Enabled2100d,
			match=>matchd2100d,
			run=>run);

	Enabled2100d <= matchd2099d;
	-- d2101d
	sted2101d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2101d,
			Enable=>Enabled2101d,
			match=>matchd2101d,
			run=>run);

	Enabled2101d <= matchd2100d;
	-- d2102d
	sted2102d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2102d,
			Enable=>Enabled2102d,
			match=>matchd2102d,
			run=>run);

	Enabled2102d <= matchd2101d;
	-- d2103d
	sted2103d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2103d,
			Enable=>Enabled2103d,
			match=>matchd2103d,
			run=>run);

	Enabled2103d <= matchd2103d OR matchd2102d;
	-- d2104d
	sted2104d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2104d,
			Enable=>Enabled2104d,
			match=>matchd2104d,
			run=>run);

	Enabled2104d <= matchd2103d;
	-- d2105d
	sted2105d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2105d,
			Enable=>Enabled2105d,
			match=>matchd2105d,
			run=>run);

	Enabled2105d <= matchd2104d;
	-- d2106d
	sted2106d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2106d,
			Enable=>Enabled2106d,
			match=>matchd2106d,
			run=>run);

	Enabled2106d <= matchd2105d;
	-- d2107d
	sted2107d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2107d,
			Enable=>Enabled2107d,
			match=>matchd2107d,
			run=>run);

	reports(109) <= matchd2107d;
	Enabled2107d <= matchd2106d;
	-- d2108d
	sted2108d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2108d,
			Enable=>Enabled2108d,
			match=>matchd2108d,
			run=>run);

	-- d2109d
	sted2109d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2109d,
			Enable=>Enabled2109d,
			match=>matchd2109d,
			run=>run);

	Enabled2109d <= matchd2108d;
	-- d2110d
	sted2110d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2110d,
			Enable=>Enabled2110d,
			match=>matchd2110d,
			run=>run);

	Enabled2110d <= matchd2109d;
	-- d2111d
	sted2111d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2111d,
			Enable=>Enabled2111d,
			match=>matchd2111d,
			run=>run);

	Enabled2111d <= matchd2110d;
	-- d2112d
	sted2112d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2112d,
			Enable=>Enabled2112d,
			match=>matchd2112d,
			run=>run);

	Enabled2112d <= matchd2111d;
	-- d2113d
	sted2113d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2113d,
			Enable=>Enabled2113d,
			match=>matchd2113d,
			run=>run);

	Enabled2113d <= matchd2112d OR matchd2113d;
	-- d2114d
	sted2114d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2114d,
			Enable=>Enabled2114d,
			match=>matchd2114d,
			run=>run);

	Enabled2114d <= matchd2113d;
	-- d2115d
	sted2115d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2115d,
			Enable=>Enabled2115d,
			match=>matchd2115d,
			run=>run);

	Enabled2115d <= matchd2114d OR matchd2115d;
	-- d2116d
	sted2116d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2116d,
			Enable=>Enabled2116d,
			match=>matchd2116d,
			run=>run);

	Enabled2116d <= matchd2115d;
	-- d2117d
	sted2117d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2117d,
			Enable=>Enabled2117d,
			match=>matchd2117d,
			run=>run);

	Enabled2117d <= matchd2116d;
	-- d2118d
	sted2118d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2118d,
			Enable=>Enabled2118d,
			match=>matchd2118d,
			run=>run);

	Enabled2118d <= matchd2117d;
	-- d2119d
	sted2119d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2119d,
			Enable=>Enabled2119d,
			match=>matchd2119d,
			run=>run);

	reports(110) <= matchd2119d;
	Enabled2119d <= matchd2118d;
	-- d2120d
	sted2120d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2120d,
			Enable=>Enabled2120d,
			match=>matchd2120d,
			run=>run);

	-- d2121d
	sted2121d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2121d,
			Enable=>Enabled2121d,
			match=>matchd2121d,
			run=>run);

	Enabled2121d <= matchd2121d OR matchd2120d;
	-- d2122d
	sted2122d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2122d,
			Enable=>Enabled2122d,
			match=>matchd2122d,
			run=>run);

	Enabled2122d <= matchd2121d;
	-- d2123d
	sted2123d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2123d,
			Enable=>Enabled2123d,
			match=>matchd2123d,
			run=>run);

	Enabled2123d <= matchd2122d;
	-- d2124d
	sted2124d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2124d,
			Enable=>Enabled2124d,
			match=>matchd2124d,
			run=>run);

	Enabled2124d <= matchd2123d;
	-- d2125d
	sted2125d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2125d,
			Enable=>Enabled2125d,
			match=>matchd2125d,
			run=>run);

	Enabled2125d <= matchd2124d;
	-- d2126d
	sted2126d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2126d,
			Enable=>Enabled2126d,
			match=>matchd2126d,
			run=>run);

	Enabled2126d <= matchd2125d;
	-- d2127d
	sted2127d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2127d,
			Enable=>Enabled2127d,
			match=>matchd2127d,
			run=>run);

	Enabled2127d <= matchd2126d;
	-- d2128d
	sted2128d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2128d,
			Enable=>Enabled2128d,
			match=>matchd2128d,
			run=>run);

	Enabled2128d <= matchd2127d;
	-- d2129d
	sted2129d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2129d,
			Enable=>Enabled2129d,
			match=>matchd2129d,
			run=>run);

	Enabled2129d <= matchd2128d;
	-- d2130d
	sted2130d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2130d,
			Enable=>Enabled2130d,
			match=>matchd2130d,
			run=>run);

	Enabled2130d <= matchd2130d OR matchd2129d;
	-- d2131d
	sted2131d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2131d,
			Enable=>Enabled2131d,
			match=>matchd2131d,
			run=>run);

	Enabled2131d <= matchd2130d;
	-- d2132d
	sted2132d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2132d,
			Enable=>Enabled2132d,
			match=>matchd2132d,
			run=>run);

	Enabled2132d <= matchd2131d;
	-- d2133d
	sted2133d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2133d,
			Enable=>Enabled2133d,
			match=>matchd2133d,
			run=>run);

	Enabled2133d <= matchd2132d;
	-- d2134d
	sted2134d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2134d,
			Enable=>Enabled2134d,
			match=>matchd2134d,
			run=>run);

	Enabled2134d <= matchd2133d;
	-- d2135d
	sted2135d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2135d,
			Enable=>Enabled2135d,
			match=>matchd2135d,
			run=>run);

	Enabled2135d <= matchd2134d;
	-- d2136d
	sted2136d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2136d,
			Enable=>Enabled2136d,
			match=>matchd2136d,
			run=>run);

	Enabled2136d <= matchd2135d OR matchd2136d;
	-- d2137d
	sted2137d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2137d,
			Enable=>Enabled2137d,
			match=>matchd2137d,
			run=>run);

	Enabled2137d <= matchd2136d;
	-- d2138d
	sted2138d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2138d,
			Enable=>Enabled2138d,
			match=>matchd2138d,
			run=>run);

	Enabled2138d <= matchd2137d;
	-- d2139d
	sted2139d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2139d,
			Enable=>Enabled2139d,
			match=>matchd2139d,
			run=>run);

	Enabled2139d <= matchd2138d;
	-- d2140d
	sted2140d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2140d,
			Enable=>Enabled2140d,
			match=>matchd2140d,
			run=>run);

	Enabled2140d <= matchd2139d;
	-- d2141d
	sted2141d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2141d,
			Enable=>Enabled2141d,
			match=>matchd2141d,
			run=>run);

	reports(111) <= matchd2141d;
	Enabled2141d <= matchd2140d;
	-- d2142d
	sted2142d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2142d,
			Enable=>Enabled2142d,
			match=>matchd2142d,
			run=>run);

	-- d2143d
	sted2143d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2143d,
			Enable=>Enabled2143d,
			match=>matchd2143d,
			run=>run);

	Enabled2143d <= matchd2142d OR matchd2143d;
	-- d2144d
	sted2144d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2144d,
			Enable=>Enabled2144d,
			match=>matchd2144d,
			run=>run);

	Enabled2144d <= matchd2143d;
	-- d2145d
	sted2145d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2145d,
			Enable=>Enabled2145d,
			match=>matchd2145d,
			run=>run);

	Enabled2145d <= matchd2144d;
	-- d2146d
	sted2146d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2146d,
			Enable=>Enabled2146d,
			match=>matchd2146d,
			run=>run);

	Enabled2146d <= matchd2145d;
	-- d2147d
	sted2147d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2147d,
			Enable=>Enabled2147d,
			match=>matchd2147d,
			run=>run);

	Enabled2147d <= matchd2146d;
	-- d2148d
	sted2148d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2148d,
			Enable=>Enabled2148d,
			match=>matchd2148d,
			run=>run);

	Enabled2148d <= matchd2147d;
	-- d2149d
	sted2149d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2149d,
			Enable=>Enabled2149d,
			match=>matchd2149d,
			run=>run);

	Enabled2149d <= matchd2149d OR matchd2148d;
	-- d2150d
	sted2150d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2150d,
			Enable=>Enabled2150d,
			match=>matchd2150d,
			run=>run);

	Enabled2150d <= matchd2149d;
	-- d2151d
	sted2151d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2151d,
			Enable=>Enabled2151d,
			match=>matchd2151d,
			run=>run);

	Enabled2151d <= matchd2150d;
	-- d2152d
	sted2152d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2152d,
			Enable=>Enabled2152d,
			match=>matchd2152d,
			run=>run);

	Enabled2152d <= matchd2151d;
	-- d2153d
	sted2153d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2153d,
			Enable=>Enabled2153d,
			match=>matchd2153d,
			run=>run);

	Enabled2153d <= matchd2152d;
	-- d2154d
	sted2154d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2154d,
			Enable=>Enabled2154d,
			match=>matchd2154d,
			run=>run);

	Enabled2154d <= matchd2153d OR matchd2154d;
	-- d2155d
	sted2155d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2155d,
			Enable=>Enabled2155d,
			match=>matchd2155d,
			run=>run);

	Enabled2155d <= matchd2154d;
	-- d2156d
	sted2156d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2156d,
			Enable=>Enabled2156d,
			match=>matchd2156d,
			run=>run);

	Enabled2156d <= matchd2155d;
	-- d2157d
	sted2157d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2157d,
			Enable=>Enabled2157d,
			match=>matchd2157d,
			run=>run);

	Enabled2157d <= matchd2156d;
	-- d2158d
	sted2158d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2158d,
			Enable=>Enabled2158d,
			match=>matchd2158d,
			run=>run);

	reports(112) <= matchd2158d;
	Enabled2158d <= matchd2157d;
	-- d2159d
	sted2159d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2159d,
			Enable=>Enabled2159d,
			match=>matchd2159d,
			run=>run);

	-- d2160d
	sted2160d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2160d,
			Enable=>Enabled2160d,
			match=>matchd2160d,
			run=>run);

	Enabled2160d <= matchd2159d OR matchd2160d;
	-- d2161d
	sted2161d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2161d,
			Enable=>Enabled2161d,
			match=>matchd2161d,
			run=>run);

	Enabled2161d <= matchd2160d;
	-- d2162d
	sted2162d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2162d,
			Enable=>Enabled2162d,
			match=>matchd2162d,
			run=>run);

	Enabled2162d <= matchd2161d;
	-- d2163d
	sted2163d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2163d,
			Enable=>Enabled2163d,
			match=>matchd2163d,
			run=>run);

	Enabled2163d <= matchd2162d;
	-- d2164d
	sted2164d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2164d,
			Enable=>Enabled2164d,
			match=>matchd2164d,
			run=>run);

	Enabled2164d <= matchd2163d;
	-- d2165d
	sted2165d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2165d,
			Enable=>Enabled2165d,
			match=>matchd2165d,
			run=>run);

	Enabled2165d <= matchd2165d OR matchd2164d;
	-- d2166d
	sted2166d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2166d,
			Enable=>Enabled2166d,
			match=>matchd2166d,
			run=>run);

	Enabled2166d <= matchd2165d;
	-- d2167d
	sted2167d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2167d,
			Enable=>Enabled2167d,
			match=>matchd2167d,
			run=>run);

	Enabled2167d <= matchd2166d;
	-- d2168d
	sted2168d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2168d,
			Enable=>Enabled2168d,
			match=>matchd2168d,
			run=>run);

	Enabled2168d <= matchd2167d;
	-- d2169d
	sted2169d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2169d,
			Enable=>Enabled2169d,
			match=>matchd2169d,
			run=>run);

	Enabled2169d <= matchd2168d;
	-- d2170d
	sted2170d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2170d,
			Enable=>Enabled2170d,
			match=>matchd2170d,
			run=>run);

	reports(113) <= matchd2170d;
	Enabled2170d <= matchd2169d;
	-- d2171d
	sted2171d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2171d,
			Enable=>Enabled2171d,
			match=>matchd2171d,
			run=>run);

	-- d2172d
	sted2172d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2172d,
			Enable=>Enabled2172d,
			match=>matchd2172d,
			run=>run);

	Enabled2172d <= matchd2172d OR matchd2171d;
	-- d2173d
	sted2173d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2173d,
			Enable=>Enabled2173d,
			match=>matchd2173d,
			run=>run);

	Enabled2173d <= matchd2172d;
	-- d2174d
	sted2174d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2174d,
			Enable=>Enabled2174d,
			match=>matchd2174d,
			run=>run);

	Enabled2174d <= matchd2173d;
	-- d2175d
	sted2175d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2175d,
			Enable=>Enabled2175d,
			match=>matchd2175d,
			run=>run);

	Enabled2175d <= matchd2174d;
	-- d2176d
	sted2176d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2176d,
			Enable=>Enabled2176d,
			match=>matchd2176d,
			run=>run);

	Enabled2176d <= matchd2175d;
	-- d2177d
	sted2177d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2177d,
			Enable=>Enabled2177d,
			match=>matchd2177d,
			run=>run);

	Enabled2177d <= matchd2176d;
	-- d2178d
	sted2178d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2178d,
			Enable=>Enabled2178d,
			match=>matchd2178d,
			run=>run);

	Enabled2178d <= matchd2177d;
	-- d2179d
	sted2179d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2179d,
			Enable=>Enabled2179d,
			match=>matchd2179d,
			run=>run);

	Enabled2179d <= matchd2178d;
	-- d2180d
	sted2180d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2180d,
			Enable=>Enabled2180d,
			match=>matchd2180d,
			run=>run);

	Enabled2180d <= matchd2179d;
	-- d2181d
	sted2181d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2181d,
			Enable=>Enabled2181d,
			match=>matchd2181d,
			run=>run);

	Enabled2181d <= matchd2181d OR matchd2180d;
	-- d2182d
	sted2182d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2182d,
			Enable=>Enabled2182d,
			match=>matchd2182d,
			run=>run);

	Enabled2182d <= matchd2181d;
	-- d2183d
	sted2183d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2183d,
			Enable=>Enabled2183d,
			match=>matchd2183d,
			run=>run);

	Enabled2183d <= matchd2182d;
	-- d2184d
	sted2184d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2184d,
			Enable=>Enabled2184d,
			match=>matchd2184d,
			run=>run);

	Enabled2184d <= matchd2183d;
	-- d2185d
	sted2185d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2185d,
			Enable=>Enabled2185d,
			match=>matchd2185d,
			run=>run);

	Enabled2185d <= matchd2184d;
	-- d2186d
	sted2186d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2186d,
			Enable=>Enabled2186d,
			match=>matchd2186d,
			run=>run);

	Enabled2186d <= matchd2185d;
	-- d2187d
	sted2187d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2187d,
			Enable=>Enabled2187d,
			match=>matchd2187d,
			run=>run);

	Enabled2187d <= matchd2187d OR matchd2186d;
	-- d2188d
	sted2188d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2188d,
			Enable=>Enabled2188d,
			match=>matchd2188d,
			run=>run);

	Enabled2188d <= matchd2187d;
	-- d2189d
	sted2189d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2189d,
			Enable=>Enabled2189d,
			match=>matchd2189d,
			run=>run);

	Enabled2189d <= matchd2188d;
	-- d2190d
	sted2190d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2190d,
			Enable=>Enabled2190d,
			match=>matchd2190d,
			run=>run);

	Enabled2190d <= matchd2189d;
	-- d2191d
	sted2191d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2191d,
			Enable=>Enabled2191d,
			match=>matchd2191d,
			run=>run);

	Enabled2191d <= matchd2190d;
	-- d2192d
	sted2192d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2192d,
			Enable=>Enabled2192d,
			match=>matchd2192d,
			run=>run);

	reports(114) <= matchd2192d;
	Enabled2192d <= matchd2191d;
	-- d2193d
	sted2193d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2193d,
			Enable=>Enabled2193d,
			match=>matchd2193d,
			run=>run);

	-- d2194d
	sted2194d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2194d,
			Enable=>Enabled2194d,
			match=>matchd2194d,
			run=>run);

	Enabled2194d <= matchd2193d;
	-- d2195d
	sted2195d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2195d,
			Enable=>Enabled2195d,
			match=>matchd2195d,
			run=>run);

	Enabled2195d <= matchd2194d;
	-- d2196d
	sted2196d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2196d,
			Enable=>Enabled2196d,
			match=>matchd2196d,
			run=>run);

	Enabled2196d <= matchd2195d;
	-- d2197d
	sted2197d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2197d,
			Enable=>Enabled2197d,
			match=>matchd2197d,
			run=>run);

	Enabled2197d <= matchd2196d;
	-- d2198d
	sted2198d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2198d,
			Enable=>Enabled2198d,
			match=>matchd2198d,
			run=>run);

	Enabled2198d <= matchd2197d;
	-- d2199d
	sted2199d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2199d,
			Enable=>Enabled2199d,
			match=>matchd2199d,
			run=>run);

	Enabled2199d <= matchd2198d;
	-- d2200d
	sted2200d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2200d,
			Enable=>Enabled2200d,
			match=>matchd2200d,
			run=>run);

	Enabled2200d <= matchd2199d OR matchd2200d;
	-- d2201d
	sted2201d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2201d,
			Enable=>Enabled2201d,
			match=>matchd2201d,
			run=>run);

	Enabled2201d <= matchd2200d;
	-- d2202d
	sted2202d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2202d,
			Enable=>Enabled2202d,
			match=>matchd2202d,
			run=>run);

	Enabled2202d <= matchd2201d OR matchd2202d;
	-- d2203d
	sted2203d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2203d,
			Enable=>Enabled2203d,
			match=>matchd2203d,
			run=>run);

	Enabled2203d <= matchd2202d;
	-- d2204d
	sted2204d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2204d,
			Enable=>Enabled2204d,
			match=>matchd2204d,
			run=>run);

	Enabled2204d <= matchd2203d;
	-- d2205d
	sted2205d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2205d,
			Enable=>Enabled2205d,
			match=>matchd2205d,
			run=>run);

	Enabled2205d <= matchd2204d;
	-- d2206d
	sted2206d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2206d,
			Enable=>Enabled2206d,
			match=>matchd2206d,
			run=>run);

	Enabled2206d <= matchd2205d;
	-- d2207d
	sted2207d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2207d,
			Enable=>Enabled2207d,
			match=>matchd2207d,
			run=>run);

	Enabled2207d <= matchd2206d OR matchd2207d;
	-- d2208d
	sted2208d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2208d,
			Enable=>Enabled2208d,
			match=>matchd2208d,
			run=>run);

	reports(115) <= matchd2208d;
	Enabled2208d <= matchd2207d;
	-- d2209d
	sted2209d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2209d,
			Enable=>Enabled2209d,
			match=>matchd2209d,
			run=>run);

	-- d2210d
	sted2210d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2210d,
			Enable=>Enabled2210d,
			match=>matchd2210d,
			run=>run);

	Enabled2210d <= matchd2209d OR matchd2210d;
	-- d2211d
	sted2211d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2211d,
			Enable=>Enabled2211d,
			match=>matchd2211d,
			run=>run);

	Enabled2211d <= matchd2210d;
	-- d2212d
	sted2212d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2212d,
			Enable=>Enabled2212d,
			match=>matchd2212d,
			run=>run);

	Enabled2212d <= matchd2211d;
	-- d2213d
	sted2213d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2213d,
			Enable=>Enabled2213d,
			match=>matchd2213d,
			run=>run);

	Enabled2213d <= matchd2212d;
	-- d2214d
	sted2214d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2214d,
			Enable=>Enabled2214d,
			match=>matchd2214d,
			run=>run);

	Enabled2214d <= matchd2213d;
	-- d2215d
	sted2215d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2215d,
			Enable=>Enabled2215d,
			match=>matchd2215d,
			run=>run);

	Enabled2215d <= matchd2215d OR matchd2214d;
	-- d2216d
	sted2216d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2216d,
			Enable=>Enabled2216d,
			match=>matchd2216d,
			run=>run);

	Enabled2216d <= matchd2215d;
	-- d2217d
	sted2217d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2217d,
			Enable=>Enabled2217d,
			match=>matchd2217d,
			run=>run);

	Enabled2217d <= matchd2216d;
	-- d2218d
	sted2218d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2218d,
			Enable=>Enabled2218d,
			match=>matchd2218d,
			run=>run);

	Enabled2218d <= matchd2217d;
	-- d2219d
	sted2219d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2219d,
			Enable=>Enabled2219d,
			match=>matchd2219d,
			run=>run);

	Enabled2219d <= matchd2218d;
	-- d2220d
	sted2220d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2220d,
			Enable=>Enabled2220d,
			match=>matchd2220d,
			run=>run);

	reports(116) <= matchd2220d;
	Enabled2220d <= matchd2219d;
	-- d2221d
	sted2221d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2221d,
			Enable=>Enabled2221d,
			match=>matchd2221d,
			run=>run);

	-- d2222d
	sted2222d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2222d,
			Enable=>Enabled2222d,
			match=>matchd2222d,
			run=>run);

	Enabled2222d <= matchd2221d;
	-- d2223d
	sted2223d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2223d,
			Enable=>Enabled2223d,
			match=>matchd2223d,
			run=>run);

	Enabled2223d <= matchd2222d;
	-- d2224d
	sted2224d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2224d,
			Enable=>Enabled2224d,
			match=>matchd2224d,
			run=>run);

	Enabled2224d <= matchd2223d;
	-- d2225d
	sted2225d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2225d,
			Enable=>Enabled2225d,
			match=>matchd2225d,
			run=>run);

	Enabled2225d <= matchd2224d;
	-- d2226d
	sted2226d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2226d,
			Enable=>Enabled2226d,
			match=>matchd2226d,
			run=>run);

	Enabled2226d <= matchd2225d;
	-- d2227d
	sted2227d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2227d,
			Enable=>Enabled2227d,
			match=>matchd2227d,
			run=>run);

	Enabled2227d <= matchd2226d;
	-- d2228d
	sted2228d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2228d,
			Enable=>Enabled2228d,
			match=>matchd2228d,
			run=>run);

	Enabled2228d <= matchd2227d;
	-- d2229d
	sted2229d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2229d,
			Enable=>Enabled2229d,
			match=>matchd2229d,
			run=>run);

	Enabled2229d <= matchd2228d;
	-- d2230d
	sted2230d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2230d,
			Enable=>Enabled2230d,
			match=>matchd2230d,
			run=>run);

	Enabled2230d <= matchd2229d;
	-- d2231d
	sted2231d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2231d,
			Enable=>Enabled2231d,
			match=>matchd2231d,
			run=>run);

	Enabled2231d <= matchd2230d;
	-- d2232d
	sted2232d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2232d,
			Enable=>Enabled2232d,
			match=>matchd2232d,
			run=>run);

	reports(117) <= matchd2232d;
	Enabled2232d <= matchd2231d;
	-- d2233d
	sted2233d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2233d,
			Enable=>Enabled2233d,
			match=>matchd2233d,
			run=>run);

	-- d2234d
	sted2234d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2234d,
			Enable=>Enabled2234d,
			match=>matchd2234d,
			run=>run);

	Enabled2234d <= matchd2233d OR matchd2234d;
	-- d2235d
	sted2235d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2235d,
			Enable=>Enabled2235d,
			match=>matchd2235d,
			run=>run);

	Enabled2235d <= matchd2234d;
	-- d2236d
	sted2236d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2236d,
			Enable=>Enabled2236d,
			match=>matchd2236d,
			run=>run);

	Enabled2236d <= matchd2235d;
	-- d2237d
	sted2237d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2237d,
			Enable=>Enabled2237d,
			match=>matchd2237d,
			run=>run);

	Enabled2237d <= matchd2236d;
	-- d2238d
	sted2238d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2238d,
			Enable=>Enabled2238d,
			match=>matchd2238d,
			run=>run);

	Enabled2238d <= matchd2237d;
	-- d2239d
	sted2239d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2239d,
			Enable=>Enabled2239d,
			match=>matchd2239d,
			run=>run);

	Enabled2239d <= matchd2239d OR matchd2238d;
	-- d2240d
	sted2240d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2240d,
			Enable=>Enabled2240d,
			match=>matchd2240d,
			run=>run);

	Enabled2240d <= matchd2239d;
	-- d2241d
	sted2241d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2241d,
			Enable=>Enabled2241d,
			match=>matchd2241d,
			run=>run);

	Enabled2241d <= matchd2240d;
	-- d2242d
	sted2242d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2242d,
			Enable=>Enabled2242d,
			match=>matchd2242d,
			run=>run);

	Enabled2242d <= matchd2241d;
	-- d2243d
	sted2243d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2243d,
			Enable=>Enabled2243d,
			match=>matchd2243d,
			run=>run);

	Enabled2243d <= matchd2242d;
	-- d2244d
	sted2244d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2244d,
			Enable=>Enabled2244d,
			match=>matchd2244d,
			run=>run);

	Enabled2244d <= matchd2243d;
	-- d2245d
	sted2245d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2245d,
			Enable=>Enabled2245d,
			match=>matchd2245d,
			run=>run);

	Enabled2245d <= matchd2244d OR matchd2245d;
	-- d2246d
	sted2246d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2246d,
			Enable=>Enabled2246d,
			match=>matchd2246d,
			run=>run);

	Enabled2246d <= matchd2245d;
	-- d2247d
	sted2247d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2247d,
			Enable=>Enabled2247d,
			match=>matchd2247d,
			run=>run);

	Enabled2247d <= matchd2246d;
	-- d2248d
	sted2248d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2248d,
			Enable=>Enabled2248d,
			match=>matchd2248d,
			run=>run);

	Enabled2248d <= matchd2247d;
	-- d2249d
	sted2249d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2249d,
			Enable=>Enabled2249d,
			match=>matchd2249d,
			run=>run);

	Enabled2249d <= matchd2248d;
	-- d2250d
	sted2250d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2250d,
			Enable=>Enabled2250d,
			match=>matchd2250d,
			run=>run);

	Enabled2250d <= matchd2249d;
	-- d2251d
	sted2251d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2251d,
			Enable=>Enabled2251d,
			match=>matchd2251d,
			run=>run);

	reports(118) <= matchd2251d;
	Enabled2251d <= matchd2250d;
	-- d2252d
	sted2252d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2252d,
			Enable=>Enabled2252d,
			match=>matchd2252d,
			run=>run);

	-- d2253d
	sted2253d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2253d,
			Enable=>Enabled2253d,
			match=>matchd2253d,
			run=>run);

	Enabled2253d <= matchd2252d OR matchd2253d;
	-- d2254d
	sted2254d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2254d,
			Enable=>Enabled2254d,
			match=>matchd2254d,
			run=>run);

	Enabled2254d <= matchd2253d;
	-- d2255d
	sted2255d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2255d,
			Enable=>Enabled2255d,
			match=>matchd2255d,
			run=>run);

	Enabled2255d <= matchd2254d;
	-- d2256d
	sted2256d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2256d,
			Enable=>Enabled2256d,
			match=>matchd2256d,
			run=>run);

	Enabled2256d <= matchd2255d;
	-- d2257d
	sted2257d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2257d,
			Enable=>Enabled2257d,
			match=>matchd2257d,
			run=>run);

	Enabled2257d <= matchd2256d;
	-- d2258d
	sted2258d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2258d,
			Enable=>Enabled2258d,
			match=>matchd2258d,
			run=>run);

	Enabled2258d <= matchd2257d OR matchd2258d;
	-- d2259d
	sted2259d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2259d,
			Enable=>Enabled2259d,
			match=>matchd2259d,
			run=>run);

	Enabled2259d <= matchd2258d;
	-- d2260d
	sted2260d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2260d,
			Enable=>Enabled2260d,
			match=>matchd2260d,
			run=>run);

	Enabled2260d <= matchd2259d;
	-- d2261d
	sted2261d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2261d,
			Enable=>Enabled2261d,
			match=>matchd2261d,
			run=>run);

	Enabled2261d <= matchd2260d;
	-- d2262d
	sted2262d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2262d,
			Enable=>Enabled2262d,
			match=>matchd2262d,
			run=>run);

	Enabled2262d <= matchd2261d;
	-- d2263d
	sted2263d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2263d,
			Enable=>Enabled2263d,
			match=>matchd2263d,
			run=>run);

	reports(119) <= matchd2263d;
	Enabled2263d <= matchd2262d;
	-- d2264d
	sted2264d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2264d,
			Enable=>Enabled2264d,
			match=>matchd2264d,
			run=>run);

	-- d2265d
	sted2265d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2265d,
			Enable=>Enabled2265d,
			match=>matchd2265d,
			run=>run);

	Enabled2265d <= matchd2264d OR matchd2265d;
	-- d2266d
	sted2266d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2266d,
			Enable=>Enabled2266d,
			match=>matchd2266d,
			run=>run);

	Enabled2266d <= matchd2265d;
	-- d2267d
	sted2267d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2267d,
			Enable=>Enabled2267d,
			match=>matchd2267d,
			run=>run);

	Enabled2267d <= matchd2266d;
	-- d2268d
	sted2268d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2268d,
			Enable=>Enabled2268d,
			match=>matchd2268d,
			run=>run);

	Enabled2268d <= matchd2267d;
	-- d2269d
	sted2269d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2269d,
			Enable=>Enabled2269d,
			match=>matchd2269d,
			run=>run);

	Enabled2269d <= matchd2268d;
	-- d2270d
	sted2270d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2270d,
			Enable=>Enabled2270d,
			match=>matchd2270d,
			run=>run);

	Enabled2270d <= matchd2269d;
	-- d2271d
	sted2271d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2271d,
			Enable=>Enabled2271d,
			match=>matchd2271d,
			run=>run);

	Enabled2271d <= matchd2270d;
	-- d2272d
	sted2272d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2272d,
			Enable=>Enabled2272d,
			match=>matchd2272d,
			run=>run);

	Enabled2272d <= matchd2271d;
	-- d2273d
	sted2273d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2273d,
			Enable=>Enabled2273d,
			match=>matchd2273d,
			run=>run);

	Enabled2273d <= matchd2272d;
	-- d2274d
	sted2274d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2274d,
			Enable=>Enabled2274d,
			match=>matchd2274d,
			run=>run);

	Enabled2274d <= matchd2273d;
	-- d2275d
	sted2275d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2275d,
			Enable=>Enabled2275d,
			match=>matchd2275d,
			run=>run);

	Enabled2275d <= matchd2274d;
	-- d2276d
	sted2276d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2276d,
			Enable=>Enabled2276d,
			match=>matchd2276d,
			run=>run);

	Enabled2276d <= matchd2275d;
	-- d2277d
	sted2277d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2277d,
			Enable=>Enabled2277d,
			match=>matchd2277d,
			run=>run);

	Enabled2277d <= matchd2276d;
	-- d2278d
	sted2278d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2278d,
			Enable=>Enabled2278d,
			match=>matchd2278d,
			run=>run);

	Enabled2278d <= matchd2277d;
	-- d2279d
	sted2279d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2279d,
			Enable=>Enabled2279d,
			match=>matchd2279d,
			run=>run);

	reports(120) <= matchd2279d;
	Enabled2279d <= matchd2278d;
	-- d2280d
	sted2280d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2280d,
			Enable=>Enabled2280d,
			match=>matchd2280d,
			run=>run);

	-- d2281d
	sted2281d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2281d,
			Enable=>Enabled2281d,
			match=>matchd2281d,
			run=>run);

	Enabled2281d <= matchd2280d;
	-- d2282d
	sted2282d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2282d,
			Enable=>Enabled2282d,
			match=>matchd2282d,
			run=>run);

	Enabled2282d <= matchd2281d;
	-- d2283d
	sted2283d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2283d,
			Enable=>Enabled2283d,
			match=>matchd2283d,
			run=>run);

	Enabled2283d <= matchd2282d;
	-- d2284d
	sted2284d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2284d,
			Enable=>Enabled2284d,
			match=>matchd2284d,
			run=>run);

	Enabled2284d <= matchd2283d;
	-- d2285d
	sted2285d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2285d,
			Enable=>Enabled2285d,
			match=>matchd2285d,
			run=>run);

	Enabled2285d <= matchd2284d OR matchd2285d;
	-- d2286d
	sted2286d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2286d,
			Enable=>Enabled2286d,
			match=>matchd2286d,
			run=>run);

	Enabled2286d <= matchd2285d;
	-- d2287d
	sted2287d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2287d,
			Enable=>Enabled2287d,
			match=>matchd2287d,
			run=>run);

	Enabled2287d <= matchd2287d OR matchd2286d;
	-- d2288d
	sted2288d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2288d,
			Enable=>Enabled2288d,
			match=>matchd2288d,
			run=>run);

	Enabled2288d <= matchd2287d;
	-- d2289d
	sted2289d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2289d,
			Enable=>Enabled2289d,
			match=>matchd2289d,
			run=>run);

	Enabled2289d <= matchd2288d;
	-- d2290d
	sted2290d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2290d,
			Enable=>Enabled2290d,
			match=>matchd2290d,
			run=>run);

	Enabled2290d <= matchd2289d;
	-- d2291d
	sted2291d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2291d,
			Enable=>Enabled2291d,
			match=>matchd2291d,
			run=>run);

	reports(121) <= matchd2291d;
	Enabled2291d <= matchd2290d;
	-- d2292d
	sted2292d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2292d,
			Enable=>Enabled2292d,
			match=>matchd2292d,
			run=>run);

	-- d2293d
	sted2293d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2293d,
			Enable=>Enabled2293d,
			match=>matchd2293d,
			run=>run);

	Enabled2293d <= matchd2292d OR matchd2293d;
	-- d2294d
	sted2294d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2294d,
			Enable=>Enabled2294d,
			match=>matchd2294d,
			run=>run);

	Enabled2294d <= matchd2293d;
	-- d2295d
	sted2295d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2295d,
			Enable=>Enabled2295d,
			match=>matchd2295d,
			run=>run);

	Enabled2295d <= matchd2295d OR matchd2294d;
	-- d2296d
	sted2296d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2296d,
			Enable=>Enabled2296d,
			match=>matchd2296d,
			run=>run);

	Enabled2296d <= matchd2295d;
	-- d2297d
	sted2297d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2297d,
			Enable=>Enabled2297d,
			match=>matchd2297d,
			run=>run);

	Enabled2297d <= matchd2296d;
	-- d2298d
	sted2298d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2298d,
			Enable=>Enabled2298d,
			match=>matchd2298d,
			run=>run);

	Enabled2298d <= matchd2297d;
	-- d2299d
	sted2299d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2299d,
			Enable=>Enabled2299d,
			match=>matchd2299d,
			run=>run);

	Enabled2299d <= matchd2298d;
	-- d2300d
	sted2300d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2300d,
			Enable=>Enabled2300d,
			match=>matchd2300d,
			run=>run);

	Enabled2300d <= matchd2300d OR matchd2299d;
	-- d2301d
	sted2301d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2301d,
			Enable=>Enabled2301d,
			match=>matchd2301d,
			run=>run);

	Enabled2301d <= matchd2300d;
	-- d2302d
	sted2302d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2302d,
			Enable=>Enabled2302d,
			match=>matchd2302d,
			run=>run);

	Enabled2302d <= matchd2302d OR matchd2301d;
	-- d2303d
	sted2303d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2303d,
			Enable=>Enabled2303d,
			match=>matchd2303d,
			run=>run);

	Enabled2303d <= matchd2302d;
	-- d2304d
	sted2304d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2304d,
			Enable=>Enabled2304d,
			match=>matchd2304d,
			run=>run);

	Enabled2304d <= matchd2303d;
	-- d2305d
	sted2305d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2305d,
			Enable=>Enabled2305d,
			match=>matchd2305d,
			run=>run);

	Enabled2305d <= matchd2304d;
	-- d2306d
	sted2306d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2306d,
			Enable=>Enabled2306d,
			match=>matchd2306d,
			run=>run);

	Enabled2306d <= matchd2305d;
	-- d2307d
	sted2307d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2307d,
			Enable=>Enabled2307d,
			match=>matchd2307d,
			run=>run);

	Enabled2307d <= matchd2306d;
	-- d2308d
	sted2308d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2308d,
			Enable=>Enabled2308d,
			match=>matchd2308d,
			run=>run);

	-- d2309d
	sted2309d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2309d,
			Enable=>Enabled2309d,
			match=>matchd2309d,
			run=>run);

	Enabled2309d <= matchd2308d;
	-- d2310d
	sted2310d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2310d,
			Enable=>Enabled2310d,
			match=>matchd2310d,
			run=>run);

	Enabled2310d <= matchd2309d;
	-- d2311d
	sted2311d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2311d,
			Enable=>Enabled2311d,
			match=>matchd2311d,
			run=>run);

	Enabled2311d <= matchd2310d;
	-- d2312d
	sted2312d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2312d,
			Enable=>Enabled2312d,
			match=>matchd2312d,
			run=>run);

	Enabled2312d <= matchd2312d OR matchd2311d;
	-- d2313d
	sted2313d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2313d,
			Enable=>Enabled2313d,
			match=>matchd2313d,
			run=>run);

	Enabled2313d <= matchd2312d;
	-- d2314d
	sted2314d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2314d,
			Enable=>Enabled2314d,
			match=>matchd2314d,
			run=>run);

	Enabled2314d <= matchd2313d OR matchd2314d;
	-- d2315d
	sted2315d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2315d,
			Enable=>Enabled2315d,
			match=>matchd2315d,
			run=>run);

	Enabled2315d <= matchd2314d;
	-- d2316d
	sted2316d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2316d,
			Enable=>Enabled2316d,
			match=>matchd2316d,
			run=>run);

	Enabled2316d <= matchd2315d OR matchd2316d;
	-- d2317d
	sted2317d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2317d,
			Enable=>Enabled2317d,
			match=>matchd2317d,
			run=>run);

	Enabled2317d <= matchd2316d;
	-- d2318d
	sted2318d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2318d,
			Enable=>Enabled2318d,
			match=>matchd2318d,
			run=>run);

	Enabled2318d <= matchd2318d OR matchd2317d;
	-- d2319d
	sted2319d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2319d,
			Enable=>Enabled2319d,
			match=>matchd2319d,
			run=>run);

	Enabled2319d <= matchd2318d;
	-- d2320d
	sted2320d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2320d,
			Enable=>Enabled2320d,
			match=>matchd2320d,
			run=>run);

	Enabled2320d <= matchd2319d;
	-- d2321d
	sted2321d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2321d,
			Enable=>Enabled2321d,
			match=>matchd2321d,
			run=>run);

	Enabled2321d <= matchd2320d;
	-- d2322d
	sted2322d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2322d,
			Enable=>Enabled2322d,
			match=>matchd2322d,
			run=>run);

	Enabled2322d <= matchd2321d;
	-- d2323d
	sted2323d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2323d,
			Enable=>Enabled2323d,
			match=>matchd2323d,
			run=>run);

	Enabled2323d <= matchd2322d;
	-- d2325d
	sted2325d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2325d,
			Enable=>Enabled2325d,
			match=>matchd2325d,
			run=>run);

	-- d2326d
	sted2326d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2326d,
			Enable=>Enabled2326d,
			match=>matchd2326d,
			run=>run);

	Enabled2326d <= matchd2326d OR matchd2325d;
	-- d2327d
	sted2327d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2327d,
			Enable=>Enabled2327d,
			match=>matchd2327d,
			run=>run);

	Enabled2327d <= matchd2326d;
	-- d2328d
	sted2328d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2328d,
			Enable=>Enabled2328d,
			match=>matchd2328d,
			run=>run);

	Enabled2328d <= matchd2327d;
	-- d2329d
	sted2329d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2329d,
			Enable=>Enabled2329d,
			match=>matchd2329d,
			run=>run);

	Enabled2329d <= matchd2328d;
	-- d2330d
	sted2330d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2330d,
			Enable=>Enabled2330d,
			match=>matchd2330d,
			run=>run);

	Enabled2330d <= matchd2329d;
	-- d2331d
	sted2331d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2331d,
			Enable=>Enabled2331d,
			match=>matchd2331d,
			run=>run);

	Enabled2331d <= matchd2330d OR matchd2331d;
	-- d2332d
	sted2332d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2332d,
			Enable=>Enabled2332d,
			match=>matchd2332d,
			run=>run);

	Enabled2332d <= matchd2331d;
	-- d2333d
	sted2333d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2333d,
			Enable=>Enabled2333d,
			match=>matchd2333d,
			run=>run);

	Enabled2333d <= matchd2332d;
	-- d2334d
	sted2334d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2334d,
			Enable=>Enabled2334d,
			match=>matchd2334d,
			run=>run);

	Enabled2334d <= matchd2333d;
	-- d2335d
	sted2335d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2335d,
			Enable=>Enabled2335d,
			match=>matchd2335d,
			run=>run);

	Enabled2335d <= matchd2334d;
	-- d2336d
	sted2336d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2336d,
			Enable=>Enabled2336d,
			match=>matchd2336d,
			run=>run);

	reports(122) <= matchd2336d;
	Enabled2336d <= matchd2335d;
	-- d2337d
	sted2337d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2337d,
			Enable=>Enabled2337d,
			match=>matchd2337d,
			run=>run);

	-- d2338d
	sted2338d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2338d,
			Enable=>Enabled2338d,
			match=>matchd2338d,
			run=>run);

	Enabled2338d <= matchd2337d;
	-- d2339d
	sted2339d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2339d,
			Enable=>Enabled2339d,
			match=>matchd2339d,
			run=>run);

	Enabled2339d <= matchd2338d;
	-- d2340d
	sted2340d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2340d,
			Enable=>Enabled2340d,
			match=>matchd2340d,
			run=>run);

	Enabled2340d <= matchd2339d;
	-- d2341d
	sted2341d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2341d,
			Enable=>Enabled2341d,
			match=>matchd2341d,
			run=>run);

	Enabled2341d <= matchd2340d;
	-- d2342d
	sted2342d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2342d,
			Enable=>Enabled2342d,
			match=>matchd2342d,
			run=>run);

	Enabled2342d <= matchd2341d;
	-- d2343d
	sted2343d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2343d,
			Enable=>Enabled2343d,
			match=>matchd2343d,
			run=>run);

	Enabled2343d <= matchd2342d;
	-- d2344d
	sted2344d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2344d,
			Enable=>Enabled2344d,
			match=>matchd2344d,
			run=>run);

	Enabled2344d <= matchd2343d;
	-- d2345d
	sted2345d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2345d,
			Enable=>Enabled2345d,
			match=>matchd2345d,
			run=>run);

	Enabled2345d <= matchd2344d;
	-- d2346d
	sted2346d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2346d,
			Enable=>Enabled2346d,
			match=>matchd2346d,
			run=>run);

	Enabled2346d <= matchd2345d;
	-- d2347d
	sted2347d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2347d,
			Enable=>Enabled2347d,
			match=>matchd2347d,
			run=>run);

	Enabled2347d <= matchd2346d;
	-- d2348d
	sted2348d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2348d,
			Enable=>Enabled2348d,
			match=>matchd2348d,
			run=>run);

	Enabled2348d <= matchd2347d OR matchd2348d;
	-- d2349d
	sted2349d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2349d,
			Enable=>Enabled2349d,
			match=>matchd2349d,
			run=>run);

	Enabled2349d <= matchd2348d;
	-- d2350d
	sted2350d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2350d,
			Enable=>Enabled2350d,
			match=>matchd2350d,
			run=>run);

	Enabled2350d <= matchd2349d;
	-- d2351d
	sted2351d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2351d,
			Enable=>Enabled2351d,
			match=>matchd2351d,
			run=>run);

	Enabled2351d <= matchd2350d;
	-- d2352d
	sted2352d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2352d,
			Enable=>Enabled2352d,
			match=>matchd2352d,
			run=>run);

	Enabled2352d <= matchd2351d;
	-- d2353d
	sted2353d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2353d,
			Enable=>Enabled2353d,
			match=>matchd2353d,
			run=>run);

	reports(123) <= matchd2353d;
	Enabled2353d <= matchd2352d;
	-- d2354d
	sted2354d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2354d,
			Enable=>Enabled2354d,
			match=>matchd2354d,
			run=>run);

	-- d2355d
	sted2355d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2355d,
			Enable=>Enabled2355d,
			match=>matchd2355d,
			run=>run);

	Enabled2355d <= matchd2354d;
	-- d2356d
	sted2356d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2356d,
			Enable=>Enabled2356d,
			match=>matchd2356d,
			run=>run);

	Enabled2356d <= matchd2355d;
	-- d2357d
	sted2357d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2357d,
			Enable=>Enabled2357d,
			match=>matchd2357d,
			run=>run);

	Enabled2357d <= matchd2356d;
	-- d2358d
	sted2358d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2358d,
			Enable=>Enabled2358d,
			match=>matchd2358d,
			run=>run);

	Enabled2358d <= matchd2357d;
	-- d2359d
	sted2359d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2359d,
			Enable=>Enabled2359d,
			match=>matchd2359d,
			run=>run);

	Enabled2359d <= matchd2358d OR matchd2359d;
	-- d2360d
	sted2360d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2360d,
			Enable=>Enabled2360d,
			match=>matchd2360d,
			run=>run);

	Enabled2360d <= matchd2359d;
	-- d2361d
	sted2361d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2361d,
			Enable=>Enabled2361d,
			match=>matchd2361d,
			run=>run);

	Enabled2361d <= matchd2361d OR matchd2360d;
	-- d2362d
	sted2362d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2362d,
			Enable=>Enabled2362d,
			match=>matchd2362d,
			run=>run);

	Enabled2362d <= matchd2361d;
	-- d2363d
	sted2363d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2363d,
			Enable=>Enabled2363d,
			match=>matchd2363d,
			run=>run);

	Enabled2363d <= matchd2362d;
	-- d2364d
	sted2364d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2364d,
			Enable=>Enabled2364d,
			match=>matchd2364d,
			run=>run);

	Enabled2364d <= matchd2363d;
	-- d2365d
	sted2365d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2365d,
			Enable=>Enabled2365d,
			match=>matchd2365d,
			run=>run);

	Enabled2365d <= matchd2364d;
	-- d2366d
	sted2366d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2366d,
			Enable=>Enabled2366d,
			match=>matchd2366d,
			run=>run);

	reports(124) <= matchd2366d;
	Enabled2366d <= matchd2365d;
	-- d2367d
	sted2367d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2367d,
			Enable=>Enabled2367d,
			match=>matchd2367d,
			run=>run);

	-- d2368d
	sted2368d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2368d,
			Enable=>Enabled2368d,
			match=>matchd2368d,
			run=>run);

	Enabled2368d <= matchd2367d OR matchd2368d;
	-- d2369d
	sted2369d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2369d,
			Enable=>Enabled2369d,
			match=>matchd2369d,
			run=>run);

	Enabled2369d <= matchd2368d;
	-- d2370d
	sted2370d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2370d,
			Enable=>Enabled2370d,
			match=>matchd2370d,
			run=>run);

	Enabled2370d <= matchd2369d OR matchd2370d;
	-- d2371d
	sted2371d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2371d,
			Enable=>Enabled2371d,
			match=>matchd2371d,
			run=>run);

	Enabled2371d <= matchd2370d;
	-- d2372d
	sted2372d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2372d,
			Enable=>Enabled2372d,
			match=>matchd2372d,
			run=>run);

	Enabled2372d <= matchd2371d;
	-- d2373d
	sted2373d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2373d,
			Enable=>Enabled2373d,
			match=>matchd2373d,
			run=>run);

	Enabled2373d <= matchd2372d;
	-- d2374d
	sted2374d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2374d,
			Enable=>Enabled2374d,
			match=>matchd2374d,
			run=>run);

	Enabled2374d <= matchd2373d;
	-- d2375d
	sted2375d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2375d,
			Enable=>Enabled2375d,
			match=>matchd2375d,
			run=>run);

	Enabled2375d <= matchd2374d OR matchd2375d;
	-- d2376d
	sted2376d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2376d,
			Enable=>Enabled2376d,
			match=>matchd2376d,
			run=>run);

	Enabled2376d <= matchd2375d;
	-- d2377d
	sted2377d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2377d,
			Enable=>Enabled2377d,
			match=>matchd2377d,
			run=>run);

	Enabled2377d <= matchd2376d OR matchd2377d;
	-- d2378d
	sted2378d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2378d,
			Enable=>Enabled2378d,
			match=>matchd2378d,
			run=>run);

	Enabled2378d <= matchd2377d;
	-- d2379d
	sted2379d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2379d,
			Enable=>Enabled2379d,
			match=>matchd2379d,
			run=>run);

	Enabled2379d <= matchd2378d;
	-- d2380d
	sted2380d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2380d,
			Enable=>Enabled2380d,
			match=>matchd2380d,
			run=>run);

	Enabled2380d <= matchd2379d;
	-- d2381d
	sted2381d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2381d,
			Enable=>Enabled2381d,
			match=>matchd2381d,
			run=>run);

	Enabled2381d <= matchd2380d;
	-- d2382d
	sted2382d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2382d,
			Enable=>Enabled2382d,
			match=>matchd2382d,
			run=>run);

	-- d2383d
	sted2383d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2383d,
			Enable=>Enabled2383d,
			match=>matchd2383d,
			run=>run);

	Enabled2383d <= matchd2382d;
	-- d2384d
	sted2384d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2384d,
			Enable=>Enabled2384d,
			match=>matchd2384d,
			run=>run);

	Enabled2384d <= matchd2383d;
	-- d2385d
	sted2385d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2385d,
			Enable=>Enabled2385d,
			match=>matchd2385d,
			run=>run);

	Enabled2385d <= matchd2384d;
	-- d2386d
	sted2386d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2386d,
			Enable=>Enabled2386d,
			match=>matchd2386d,
			run=>run);

	Enabled2386d <= matchd2385d OR matchd2386d;
	-- d2387d
	sted2387d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2387d,
			Enable=>Enabled2387d,
			match=>matchd2387d,
			run=>run);

	Enabled2387d <= matchd2386d;
	-- d2388d
	sted2388d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2388d,
			Enable=>Enabled2388d,
			match=>matchd2388d,
			run=>run);

	Enabled2388d <= matchd2387d OR matchd2388d;
	-- d2389d
	sted2389d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2389d,
			Enable=>Enabled2389d,
			match=>matchd2389d,
			run=>run);

	Enabled2389d <= matchd2388d;
	-- d2390d
	sted2390d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2390d,
			Enable=>Enabled2390d,
			match=>matchd2390d,
			run=>run);

	Enabled2390d <= matchd2390d OR matchd2389d;
	-- d2391d
	sted2391d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2391d,
			Enable=>Enabled2391d,
			match=>matchd2391d,
			run=>run);

	Enabled2391d <= matchd2390d;
	-- d2392d
	sted2392d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2392d,
			Enable=>Enabled2392d,
			match=>matchd2392d,
			run=>run);

	Enabled2392d <= matchd2391d OR matchd2392d;
	-- d2393d
	sted2393d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2393d,
			Enable=>Enabled2393d,
			match=>matchd2393d,
			run=>run);

	Enabled2393d <= matchd2392d;
	-- d2394d
	sted2394d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2394d,
			Enable=>Enabled2394d,
			match=>matchd2394d,
			run=>run);

	Enabled2394d <= matchd2393d;
	-- d2395d
	sted2395d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2395d,
			Enable=>Enabled2395d,
			match=>matchd2395d,
			run=>run);

	Enabled2395d <= matchd2394d;
	-- d2396d
	sted2396d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2396d,
			Enable=>Enabled2396d,
			match=>matchd2396d,
			run=>run);

	Enabled2396d <= matchd2395d;
	-- d2398d
	sted2398d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2398d,
			Enable=>Enabled2398d,
			match=>matchd2398d,
			run=>run);

	-- d2399d
	sted2399d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2399d,
			Enable=>Enabled2399d,
			match=>matchd2399d,
			run=>run);

	Enabled2399d <= matchd2398d OR matchd2399d;
	-- d2400d
	sted2400d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2400d,
			Enable=>Enabled2400d,
			match=>matchd2400d,
			run=>run);

	Enabled2400d <= matchd2399d;
	-- d2401d
	sted2401d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2401d,
			Enable=>Enabled2401d,
			match=>matchd2401d,
			run=>run);

	Enabled2401d <= matchd2400d;
	-- d2402d
	sted2402d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2402d,
			Enable=>Enabled2402d,
			match=>matchd2402d,
			run=>run);

	Enabled2402d <= matchd2401d;
	-- d2403d
	sted2403d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2403d,
			Enable=>Enabled2403d,
			match=>matchd2403d,
			run=>run);

	Enabled2403d <= matchd2402d;
	-- d2404d
	sted2404d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2404d,
			Enable=>Enabled2404d,
			match=>matchd2404d,
			run=>run);

	Enabled2404d <= matchd2404d OR matchd2403d;
	-- d2405d
	sted2405d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2405d,
			Enable=>Enabled2405d,
			match=>matchd2405d,
			run=>run);

	Enabled2405d <= matchd2404d;
	-- d2406d
	sted2406d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2406d,
			Enable=>Enabled2406d,
			match=>matchd2406d,
			run=>run);

	Enabled2406d <= matchd2405d;
	-- d2407d
	sted2407d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2407d,
			Enable=>Enabled2407d,
			match=>matchd2407d,
			run=>run);

	Enabled2407d <= matchd2406d;
	-- d2408d
	sted2408d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2408d,
			Enable=>Enabled2408d,
			match=>matchd2408d,
			run=>run);

	Enabled2408d <= matchd2407d;
	-- d2409d
	sted2409d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2409d,
			Enable=>Enabled2409d,
			match=>matchd2409d,
			run=>run);

	reports(125) <= matchd2409d;
	Enabled2409d <= matchd2408d;
	-- d2410d
	sted2410d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2410d,
			Enable=>Enabled2410d,
			match=>matchd2410d,
			run=>run);

	-- d2411d
	sted2411d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2411d,
			Enable=>Enabled2411d,
			match=>matchd2411d,
			run=>run);

	Enabled2411d <= matchd2411d OR matchd2410d;
	-- d2412d
	sted2412d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2412d,
			Enable=>Enabled2412d,
			match=>matchd2412d,
			run=>run);

	Enabled2412d <= matchd2411d;
	-- d2413d
	sted2413d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2413d,
			Enable=>Enabled2413d,
			match=>matchd2413d,
			run=>run);

	Enabled2413d <= matchd2412d;
	-- d2414d
	sted2414d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2414d,
			Enable=>Enabled2414d,
			match=>matchd2414d,
			run=>run);

	Enabled2414d <= matchd2413d;
	-- d2415d
	sted2415d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2415d,
			Enable=>Enabled2415d,
			match=>matchd2415d,
			run=>run);

	Enabled2415d <= matchd2414d;
	-- d2416d
	sted2416d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2416d,
			Enable=>Enabled2416d,
			match=>matchd2416d,
			run=>run);

	Enabled2416d <= matchd2415d OR matchd2416d;
	-- d2417d
	sted2417d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2417d,
			Enable=>Enabled2417d,
			match=>matchd2417d,
			run=>run);

	Enabled2417d <= matchd2416d;
	-- d2418d
	sted2418d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2418d,
			Enable=>Enabled2418d,
			match=>matchd2418d,
			run=>run);

	Enabled2418d <= matchd2417d;
	-- d2419d
	sted2419d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2419d,
			Enable=>Enabled2419d,
			match=>matchd2419d,
			run=>run);

	Enabled2419d <= matchd2418d;
	-- d2420d
	sted2420d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2420d,
			Enable=>Enabled2420d,
			match=>matchd2420d,
			run=>run);

	reports(126) <= matchd2420d;
	Enabled2420d <= matchd2419d;
	-- d2421d
	sted2421d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2421d,
			Enable=>Enabled2421d,
			match=>matchd2421d,
			run=>run);

	-- d2422d
	sted2422d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2422d,
			Enable=>Enabled2422d,
			match=>matchd2422d,
			run=>run);

	Enabled2422d <= matchd2421d OR matchd2422d;
	-- d2423d
	sted2423d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2423d,
			Enable=>Enabled2423d,
			match=>matchd2423d,
			run=>run);

	Enabled2423d <= matchd2422d;
	-- d2424d
	sted2424d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2424d,
			Enable=>Enabled2424d,
			match=>matchd2424d,
			run=>run);

	Enabled2424d <= matchd2423d;
	-- d2425d
	sted2425d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2425d,
			Enable=>Enabled2425d,
			match=>matchd2425d,
			run=>run);

	Enabled2425d <= matchd2424d;
	-- d2426d
	sted2426d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2426d,
			Enable=>Enabled2426d,
			match=>matchd2426d,
			run=>run);

	Enabled2426d <= matchd2425d;
	-- d2427d
	sted2427d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2427d,
			Enable=>Enabled2427d,
			match=>matchd2427d,
			run=>run);

	Enabled2427d <= matchd2426d;
	-- d2428d
	sted2428d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2428d,
			Enable=>Enabled2428d,
			match=>matchd2428d,
			run=>run);

	Enabled2428d <= matchd2428d OR matchd2427d;
	-- d2429d
	sted2429d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2429d,
			Enable=>Enabled2429d,
			match=>matchd2429d,
			run=>run);

	Enabled2429d <= matchd2428d;
	-- d2430d
	sted2430d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2430d,
			Enable=>Enabled2430d,
			match=>matchd2430d,
			run=>run);

	Enabled2430d <= matchd2429d;
	-- d2431d
	sted2431d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2431d,
			Enable=>Enabled2431d,
			match=>matchd2431d,
			run=>run);

	Enabled2431d <= matchd2430d;
	-- d2432d
	sted2432d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2432d,
			Enable=>Enabled2432d,
			match=>matchd2432d,
			run=>run);

	Enabled2432d <= matchd2431d;
	-- d2433d
	sted2433d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2433d,
			Enable=>Enabled2433d,
			match=>matchd2433d,
			run=>run);

	Enabled2433d <= matchd2433d OR matchd2432d;
	-- d2434d
	sted2434d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2434d,
			Enable=>Enabled2434d,
			match=>matchd2434d,
			run=>run);

	Enabled2434d <= matchd2433d;
	-- d2435d
	sted2435d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2435d,
			Enable=>Enabled2435d,
			match=>matchd2435d,
			run=>run);

	Enabled2435d <= matchd2434d;
	-- d2436d
	sted2436d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2436d,
			Enable=>Enabled2436d,
			match=>matchd2436d,
			run=>run);

	reports(127) <= matchd2436d;
	Enabled2436d <= matchd2435d;
	-- d2437d
	sted2437d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2437d,
			Enable=>Enabled2437d,
			match=>matchd2437d,
			run=>run);

	-- d2438d
	sted2438d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2438d,
			Enable=>Enabled2438d,
			match=>matchd2438d,
			run=>run);

	Enabled2438d <= matchd2437d;
	-- d2439d
	sted2439d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2439d,
			Enable=>Enabled2439d,
			match=>matchd2439d,
			run=>run);

	Enabled2439d <= matchd2438d;
	-- d2440d
	sted2440d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2440d,
			Enable=>Enabled2440d,
			match=>matchd2440d,
			run=>run);

	Enabled2440d <= matchd2439d;
	-- d2441d
	sted2441d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2441d,
			Enable=>Enabled2441d,
			match=>matchd2441d,
			run=>run);

	Enabled2441d <= matchd2440d;
	-- d2442d
	sted2442d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2442d,
			Enable=>Enabled2442d,
			match=>matchd2442d,
			run=>run);

	Enabled2442d <= matchd2441d;
	-- d2443d
	sted2443d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2443d,
			Enable=>Enabled2443d,
			match=>matchd2443d,
			run=>run);

	Enabled2443d <= matchd2442d;
	-- d2444d
	sted2444d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2444d,
			Enable=>Enabled2444d,
			match=>matchd2444d,
			run=>run);

	Enabled2444d <= matchd2443d;
	-- d2445d
	sted2445d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2445d,
			Enable=>Enabled2445d,
			match=>matchd2445d,
			run=>run);

	reports(128) <= matchd2445d;
	Enabled2445d <= matchd2444d;
	-- d2446d
	sted2446d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2446d,
			Enable=>Enabled2446d,
			match=>matchd2446d,
			run=>run);

	-- d2447d
	sted2447d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2447d,
			Enable=>Enabled2447d,
			match=>matchd2447d,
			run=>run);

	Enabled2447d <= matchd2446d OR matchd2447d;
	-- d2448d
	sted2448d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2448d,
			Enable=>Enabled2448d,
			match=>matchd2448d,
			run=>run);

	Enabled2448d <= matchd2447d;
	-- d2449d
	sted2449d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2449d,
			Enable=>Enabled2449d,
			match=>matchd2449d,
			run=>run);

	Enabled2449d <= matchd2448d;
	-- d2450d
	sted2450d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2450d,
			Enable=>Enabled2450d,
			match=>matchd2450d,
			run=>run);

	Enabled2450d <= matchd2449d;
	-- d2451d
	sted2451d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2451d,
			Enable=>Enabled2451d,
			match=>matchd2451d,
			run=>run);

	Enabled2451d <= matchd2450d;
	-- d2452d
	sted2452d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2452d,
			Enable=>Enabled2452d,
			match=>matchd2452d,
			run=>run);

	Enabled2452d <= matchd2451d;
	-- d2453d
	sted2453d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2453d,
			Enable=>Enabled2453d,
			match=>matchd2453d,
			run=>run);

	Enabled2453d <= matchd2452d;
	-- d2454d
	sted2454d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2454d,
			Enable=>Enabled2454d,
			match=>matchd2454d,
			run=>run);

	Enabled2454d <= matchd2453d;
	-- d2455d
	sted2455d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2455d,
			Enable=>Enabled2455d,
			match=>matchd2455d,
			run=>run);

	Enabled2455d <= matchd2454d;
	-- d2456d
	sted2456d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2456d,
			Enable=>Enabled2456d,
			match=>matchd2456d,
			run=>run);

	Enabled2456d <= matchd2455d;
	-- d2457d
	sted2457d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2457d,
			Enable=>Enabled2457d,
			match=>matchd2457d,
			run=>run);

	Enabled2457d <= matchd2456d;
	-- d2458d
	sted2458d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2458d,
			Enable=>Enabled2458d,
			match=>matchd2458d,
			run=>run);

	Enabled2458d <= matchd2457d;
	-- d2459d
	sted2459d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2459d,
			Enable=>Enabled2459d,
			match=>matchd2459d,
			run=>run);

	Enabled2459d <= matchd2458d;
	-- d2460d
	sted2460d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2460d,
			Enable=>Enabled2460d,
			match=>matchd2460d,
			run=>run);

	reports(129) <= matchd2460d;
	Enabled2460d <= matchd2459d;
	-- d2461d
	sted2461d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2461d,
			Enable=>Enabled2461d,
			match=>matchd2461d,
			run=>run);

	-- d2462d
	sted2462d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2462d,
			Enable=>Enabled2462d,
			match=>matchd2462d,
			run=>run);

	Enabled2462d <= matchd2461d OR matchd2462d;
	-- d2463d
	sted2463d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2463d,
			Enable=>Enabled2463d,
			match=>matchd2463d,
			run=>run);

	Enabled2463d <= matchd2462d;
	-- d2464d
	sted2464d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2464d,
			Enable=>Enabled2464d,
			match=>matchd2464d,
			run=>run);

	Enabled2464d <= matchd2463d;
	-- d2465d
	sted2465d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2465d,
			Enable=>Enabled2465d,
			match=>matchd2465d,
			run=>run);

	Enabled2465d <= matchd2464d;
	-- d2466d
	sted2466d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2466d,
			Enable=>Enabled2466d,
			match=>matchd2466d,
			run=>run);

	Enabled2466d <= matchd2465d;
	-- d2467d
	sted2467d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2467d,
			Enable=>Enabled2467d,
			match=>matchd2467d,
			run=>run);

	Enabled2467d <= matchd2466d OR matchd2467d;
	-- d2468d
	sted2468d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2468d,
			Enable=>Enabled2468d,
			match=>matchd2468d,
			run=>run);

	Enabled2468d <= matchd2467d;
	-- d2469d
	sted2469d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2469d,
			Enable=>Enabled2469d,
			match=>matchd2469d,
			run=>run);

	Enabled2469d <= matchd2468d;
	-- d2470d
	sted2470d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2470d,
			Enable=>Enabled2470d,
			match=>matchd2470d,
			run=>run);

	Enabled2470d <= matchd2469d;
	-- d2471d
	sted2471d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2471d,
			Enable=>Enabled2471d,
			match=>matchd2471d,
			run=>run);

	Enabled2471d <= matchd2470d;
	-- d2472d
	sted2472d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2472d,
			Enable=>Enabled2472d,
			match=>matchd2472d,
			run=>run);

	reports(130) <= matchd2472d;
	Enabled2472d <= matchd2471d;
	-- d2473d
	sted2473d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2473d,
			Enable=>Enabled2473d,
			match=>matchd2473d,
			run=>run);

	-- d2474d
	sted2474d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2474d,
			Enable=>Enabled2474d,
			match=>matchd2474d,
			run=>run);

	Enabled2474d <= matchd2474d OR matchd2473d;
	-- d2475d
	sted2475d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2475d,
			Enable=>Enabled2475d,
			match=>matchd2475d,
			run=>run);

	Enabled2475d <= matchd2474d;
	-- d2476d
	sted2476d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2476d,
			Enable=>Enabled2476d,
			match=>matchd2476d,
			run=>run);

	Enabled2476d <= matchd2475d;
	-- d2477d
	sted2477d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2477d,
			Enable=>Enabled2477d,
			match=>matchd2477d,
			run=>run);

	Enabled2477d <= matchd2476d;
	-- d2478d
	sted2478d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2478d,
			Enable=>Enabled2478d,
			match=>matchd2478d,
			run=>run);

	Enabled2478d <= matchd2477d;
	-- d2479d
	sted2479d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2479d,
			Enable=>Enabled2479d,
			match=>matchd2479d,
			run=>run);

	Enabled2479d <= matchd2479d OR matchd2478d;
	-- d2480d
	sted2480d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2480d,
			Enable=>Enabled2480d,
			match=>matchd2480d,
			run=>run);

	Enabled2480d <= matchd2479d;
	-- d2481d
	sted2481d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2481d,
			Enable=>Enabled2481d,
			match=>matchd2481d,
			run=>run);

	Enabled2481d <= matchd2480d;
	-- d2482d
	sted2482d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2482d,
			Enable=>Enabled2482d,
			match=>matchd2482d,
			run=>run);

	Enabled2482d <= matchd2481d;
	-- d2483d
	sted2483d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2483d,
			Enable=>Enabled2483d,
			match=>matchd2483d,
			run=>run);

	reports(131) <= matchd2483d;
	Enabled2483d <= matchd2482d;
	-- d2484d
	sted2484d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2484d,
			Enable=>Enabled2484d,
			match=>matchd2484d,
			run=>run);

	-- d2485d
	sted2485d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2485d,
			Enable=>Enabled2485d,
			match=>matchd2485d,
			run=>run);

	Enabled2485d <= matchd2484d OR matchd2485d;
	-- d2486d
	sted2486d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2486d,
			Enable=>Enabled2486d,
			match=>matchd2486d,
			run=>run);

	Enabled2486d <= matchd2485d;
	-- d2487d
	sted2487d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2487d,
			Enable=>Enabled2487d,
			match=>matchd2487d,
			run=>run);

	Enabled2487d <= matchd2486d;
	-- d2488d
	sted2488d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2488d,
			Enable=>Enabled2488d,
			match=>matchd2488d,
			run=>run);

	Enabled2488d <= matchd2487d;
	-- d2489d
	sted2489d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2489d,
			Enable=>Enabled2489d,
			match=>matchd2489d,
			run=>run);

	Enabled2489d <= matchd2488d;
	-- d2490d
	sted2490d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2490d,
			Enable=>Enabled2490d,
			match=>matchd2490d,
			run=>run);

	Enabled2490d <= matchd2490d OR matchd2489d;
	-- d2491d
	sted2491d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2491d,
			Enable=>Enabled2491d,
			match=>matchd2491d,
			run=>run);

	Enabled2491d <= matchd2490d;
	-- d2492d
	sted2492d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2492d,
			Enable=>Enabled2492d,
			match=>matchd2492d,
			run=>run);

	Enabled2492d <= matchd2491d;
	-- d2493d
	sted2493d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2493d,
			Enable=>Enabled2493d,
			match=>matchd2493d,
			run=>run);

	Enabled2493d <= matchd2492d;
	-- d2494d
	sted2494d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2494d,
			Enable=>Enabled2494d,
			match=>matchd2494d,
			run=>run);

	Enabled2494d <= matchd2493d;
	-- d2495d
	sted2495d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2495d,
			Enable=>Enabled2495d,
			match=>matchd2495d,
			run=>run);

	Enabled2495d <= matchd2495d OR matchd2494d;
	-- d2496d
	sted2496d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2496d,
			Enable=>Enabled2496d,
			match=>matchd2496d,
			run=>run);

	Enabled2496d <= matchd2495d;
	-- d2497d
	sted2497d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2497d,
			Enable=>Enabled2497d,
			match=>matchd2497d,
			run=>run);

	Enabled2497d <= matchd2496d;
	-- d2498d
	sted2498d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2498d,
			Enable=>Enabled2498d,
			match=>matchd2498d,
			run=>run);

	Enabled2498d <= matchd2497d;
	-- d2499d
	sted2499d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2499d,
			Enable=>Enabled2499d,
			match=>matchd2499d,
			run=>run);

	reports(132) <= matchd2499d;
	Enabled2499d <= matchd2498d;
	-- d2500d
	sted2500d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2500d,
			Enable=>Enabled2500d,
			match=>matchd2500d,
			run=>run);

	-- d2501d
	sted2501d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2501d,
			Enable=>Enabled2501d,
			match=>matchd2501d,
			run=>run);

	Enabled2501d <= matchd2501d OR matchd2500d;
	-- d2502d
	sted2502d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2502d,
			Enable=>Enabled2502d,
			match=>matchd2502d,
			run=>run);

	Enabled2502d <= matchd2501d;
	-- d2503d
	sted2503d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2503d,
			Enable=>Enabled2503d,
			match=>matchd2503d,
			run=>run);

	Enabled2503d <= matchd2502d;
	-- d2504d
	sted2504d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2504d,
			Enable=>Enabled2504d,
			match=>matchd2504d,
			run=>run);

	Enabled2504d <= matchd2503d;
	-- d2505d
	sted2505d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2505d,
			Enable=>Enabled2505d,
			match=>matchd2505d,
			run=>run);

	Enabled2505d <= matchd2504d;
	-- d2506d
	sted2506d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2506d,
			Enable=>Enabled2506d,
			match=>matchd2506d,
			run=>run);

	Enabled2506d <= matchd2505d;
	-- d2507d
	sted2507d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2507d,
			Enable=>Enabled2507d,
			match=>matchd2507d,
			run=>run);

	Enabled2507d <= matchd2506d;
	-- d2508d
	sted2508d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2508d,
			Enable=>Enabled2508d,
			match=>matchd2508d,
			run=>run);

	Enabled2508d <= matchd2507d;
	-- d2509d
	sted2509d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2509d,
			Enable=>Enabled2509d,
			match=>matchd2509d,
			run=>run);

	Enabled2509d <= matchd2508d;
	-- d2510d
	sted2510d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2510d,
			Enable=>Enabled2510d,
			match=>matchd2510d,
			run=>run);

	Enabled2510d <= matchd2509d OR matchd2510d;
	-- d2511d
	sted2511d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2511d,
			Enable=>Enabled2511d,
			match=>matchd2511d,
			run=>run);

	Enabled2511d <= matchd2510d;
	-- d2512d
	sted2512d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2512d,
			Enable=>Enabled2512d,
			match=>matchd2512d,
			run=>run);

	Enabled2512d <= matchd2511d;
	-- d2513d
	sted2513d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2513d,
			Enable=>Enabled2513d,
			match=>matchd2513d,
			run=>run);

	Enabled2513d <= matchd2512d;
	-- d2514d
	sted2514d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2514d,
			Enable=>Enabled2514d,
			match=>matchd2514d,
			run=>run);

	Enabled2514d <= matchd2513d;
	-- d2515d
	sted2515d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2515d,
			Enable=>Enabled2515d,
			match=>matchd2515d,
			run=>run);

	Enabled2515d <= matchd2514d;
	-- d2516d
	sted2516d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2516d,
			Enable=>Enabled2516d,
			match=>matchd2516d,
			run=>run);

	Enabled2516d <= matchd2516d OR matchd2515d;
	-- d2517d
	sted2517d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2517d,
			Enable=>Enabled2517d,
			match=>matchd2517d,
			run=>run);

	Enabled2517d <= matchd2516d;
	-- d2518d
	sted2518d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2518d,
			Enable=>Enabled2518d,
			match=>matchd2518d,
			run=>run);

	Enabled2518d <= matchd2517d;
	-- d2519d
	sted2519d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2519d,
			Enable=>Enabled2519d,
			match=>matchd2519d,
			run=>run);

	Enabled2519d <= matchd2518d;
	-- d2520d
	sted2520d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2520d,
			Enable=>Enabled2520d,
			match=>matchd2520d,
			run=>run);

	reports(133) <= matchd2520d;
	Enabled2520d <= matchd2519d;
	-- d2521d
	sted2521d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2521d,
			Enable=>Enabled2521d,
			match=>matchd2521d,
			run=>run);

	-- d2522d
	sted2522d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2522d,
			Enable=>Enabled2522d,
			match=>matchd2522d,
			run=>run);

	Enabled2522d <= matchd2521d OR matchd2522d;
	-- d2523d
	sted2523d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2523d,
			Enable=>Enabled2523d,
			match=>matchd2523d,
			run=>run);

	Enabled2523d <= matchd2522d;
	-- d2524d
	sted2524d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2524d,
			Enable=>Enabled2524d,
			match=>matchd2524d,
			run=>run);

	Enabled2524d <= matchd2523d;
	-- d2525d
	sted2525d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2525d,
			Enable=>Enabled2525d,
			match=>matchd2525d,
			run=>run);

	Enabled2525d <= matchd2524d;
	-- d2526d
	sted2526d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2526d,
			Enable=>Enabled2526d,
			match=>matchd2526d,
			run=>run);

	Enabled2526d <= matchd2525d;
	-- d2527d
	sted2527d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2527d,
			Enable=>Enabled2527d,
			match=>matchd2527d,
			run=>run);

	Enabled2527d <= matchd2527d OR matchd2526d;
	-- d2528d
	sted2528d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2528d,
			Enable=>Enabled2528d,
			match=>matchd2528d,
			run=>run);

	Enabled2528d <= matchd2527d;
	-- d2529d
	sted2529d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2529d,
			Enable=>Enabled2529d,
			match=>matchd2529d,
			run=>run);

	Enabled2529d <= matchd2528d;
	-- d2530d
	sted2530d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2530d,
			Enable=>Enabled2530d,
			match=>matchd2530d,
			run=>run);

	Enabled2530d <= matchd2529d;
	-- d2531d
	sted2531d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2531d,
			Enable=>Enabled2531d,
			match=>matchd2531d,
			run=>run);

	Enabled2531d <= matchd2530d;
	-- d2532d
	sted2532d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2532d,
			Enable=>Enabled2532d,
			match=>matchd2532d,
			run=>run);

	reports(134) <= matchd2532d;
	Enabled2532d <= matchd2531d;
	-- d2533d
	sted2533d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2533d,
			Enable=>Enabled2533d,
			match=>matchd2533d,
			run=>run);

	-- d2534d
	sted2534d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2534d,
			Enable=>Enabled2534d,
			match=>matchd2534d,
			run=>run);

	Enabled2534d <= matchd2533d OR matchd2534d;
	-- d2535d
	sted2535d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2535d,
			Enable=>Enabled2535d,
			match=>matchd2535d,
			run=>run);

	Enabled2535d <= matchd2534d;
	-- d2536d
	sted2536d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2536d,
			Enable=>Enabled2536d,
			match=>matchd2536d,
			run=>run);

	Enabled2536d <= matchd2535d;
	-- d2537d
	sted2537d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2537d,
			Enable=>Enabled2537d,
			match=>matchd2537d,
			run=>run);

	Enabled2537d <= matchd2536d;
	-- d2538d
	sted2538d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2538d,
			Enable=>Enabled2538d,
			match=>matchd2538d,
			run=>run);

	Enabled2538d <= matchd2537d;
	-- d2539d
	sted2539d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2539d,
			Enable=>Enabled2539d,
			match=>matchd2539d,
			run=>run);

	Enabled2539d <= matchd2539d OR matchd2538d;
	-- d2540d
	sted2540d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2540d,
			Enable=>Enabled2540d,
			match=>matchd2540d,
			run=>run);

	Enabled2540d <= matchd2539d;
	-- d2541d
	sted2541d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2541d,
			Enable=>Enabled2541d,
			match=>matchd2541d,
			run=>run);

	Enabled2541d <= matchd2540d;
	-- d2542d
	sted2542d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2542d,
			Enable=>Enabled2542d,
			match=>matchd2542d,
			run=>run);

	Enabled2542d <= matchd2541d;
	-- d2543d
	sted2543d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2543d,
			Enable=>Enabled2543d,
			match=>matchd2543d,
			run=>run);

	Enabled2543d <= matchd2542d;
	-- d2544d
	sted2544d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2544d,
			Enable=>Enabled2544d,
			match=>matchd2544d,
			run=>run);

	reports(135) <= matchd2544d;
	Enabled2544d <= matchd2543d;
	-- d2545d
	sted2545d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2545d,
			Enable=>Enabled2545d,
			match=>matchd2545d,
			run=>run);

	-- d2546d
	sted2546d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2546d,
			Enable=>Enabled2546d,
			match=>matchd2546d,
			run=>run);

	Enabled2546d <= matchd2545d OR matchd2546d;
	-- d2547d
	sted2547d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2547d,
			Enable=>Enabled2547d,
			match=>matchd2547d,
			run=>run);

	Enabled2547d <= matchd2546d;
	-- d2548d
	sted2548d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2548d,
			Enable=>Enabled2548d,
			match=>matchd2548d,
			run=>run);

	Enabled2548d <= matchd2547d;
	-- d2549d
	sted2549d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2549d,
			Enable=>Enabled2549d,
			match=>matchd2549d,
			run=>run);

	Enabled2549d <= matchd2548d;
	-- d2550d
	sted2550d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2550d,
			Enable=>Enabled2550d,
			match=>matchd2550d,
			run=>run);

	Enabled2550d <= matchd2549d;
	-- d2551d
	sted2551d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2551d,
			Enable=>Enabled2551d,
			match=>matchd2551d,
			run=>run);

	Enabled2551d <= matchd2551d OR matchd2550d;
	-- d2552d
	sted2552d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2552d,
			Enable=>Enabled2552d,
			match=>matchd2552d,
			run=>run);

	Enabled2552d <= matchd2551d;
	-- d2553d
	sted2553d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2553d,
			Enable=>Enabled2553d,
			match=>matchd2553d,
			run=>run);

	Enabled2553d <= matchd2552d;
	-- d2554d
	sted2554d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2554d,
			Enable=>Enabled2554d,
			match=>matchd2554d,
			run=>run);

	Enabled2554d <= matchd2553d;
	-- d2555d
	sted2555d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2555d,
			Enable=>Enabled2555d,
			match=>matchd2555d,
			run=>run);

	Enabled2555d <= matchd2554d;
	-- d2556d
	sted2556d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2556d,
			Enable=>Enabled2556d,
			match=>matchd2556d,
			run=>run);

	Enabled2556d <= matchd2555d;
	-- d2557d
	sted2557d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2557d,
			Enable=>Enabled2557d,
			match=>matchd2557d,
			run=>run);

	Enabled2557d <= matchd2557d OR matchd2556d;
	-- d2558d
	sted2558d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2558d,
			Enable=>Enabled2558d,
			match=>matchd2558d,
			run=>run);

	Enabled2558d <= matchd2557d;
	-- d2559d
	sted2559d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2559d,
			Enable=>Enabled2559d,
			match=>matchd2559d,
			run=>run);

	Enabled2559d <= matchd2558d;
	-- d2560d
	sted2560d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2560d,
			Enable=>Enabled2560d,
			match=>matchd2560d,
			run=>run);

	Enabled2560d <= matchd2559d;
	-- d2561d
	sted2561d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2561d,
			Enable=>Enabled2561d,
			match=>matchd2561d,
			run=>run);

	reports(136) <= matchd2561d;
	Enabled2561d <= matchd2560d;
	-- d2562d
	sted2562d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2562d,
			Enable=>Enabled2562d,
			match=>matchd2562d,
			run=>run);

	-- d2563d
	sted2563d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2563d,
			Enable=>Enabled2563d,
			match=>matchd2563d,
			run=>run);

	Enabled2563d <= matchd2562d;
	-- d2564d
	sted2564d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2564d,
			Enable=>Enabled2564d,
			match=>matchd2564d,
			run=>run);

	Enabled2564d <= matchd2563d;
	-- d2565d
	sted2565d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2565d,
			Enable=>Enabled2565d,
			match=>matchd2565d,
			run=>run);

	Enabled2565d <= matchd2564d;
	-- d2566d
	sted2566d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2566d,
			Enable=>Enabled2566d,
			match=>matchd2566d,
			run=>run);

	Enabled2566d <= matchd2566d OR matchd2565d;
	-- d2567d
	sted2567d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2567d,
			Enable=>Enabled2567d,
			match=>matchd2567d,
			run=>run);

	Enabled2567d <= matchd2566d;
	-- d2568d
	sted2568d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2568d,
			Enable=>Enabled2568d,
			match=>matchd2568d,
			run=>run);

	Enabled2568d <= matchd2567d OR matchd2568d;
	-- d2569d
	sted2569d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2569d,
			Enable=>Enabled2569d,
			match=>matchd2569d,
			run=>run);

	Enabled2569d <= matchd2568d;
	-- d2570d
	sted2570d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2570d,
			Enable=>Enabled2570d,
			match=>matchd2570d,
			run=>run);

	Enabled2570d <= matchd2569d;
	-- d2571d
	sted2571d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2571d,
			Enable=>Enabled2571d,
			match=>matchd2571d,
			run=>run);

	Enabled2571d <= matchd2570d;
	-- d2572d
	sted2572d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2572d,
			Enable=>Enabled2572d,
			match=>matchd2572d,
			run=>run);

	reports(137) <= matchd2572d;
	Enabled2572d <= matchd2571d;
	-- d2573d
	sted2573d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2573d,
			Enable=>Enabled2573d,
			match=>matchd2573d,
			run=>run);

	-- d2574d
	sted2574d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2574d,
			Enable=>Enabled2574d,
			match=>matchd2574d,
			run=>run);

	Enabled2574d <= matchd2573d OR matchd2574d;
	-- d2575d
	sted2575d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2575d,
			Enable=>Enabled2575d,
			match=>matchd2575d,
			run=>run);

	Enabled2575d <= matchd2574d;
	-- d2576d
	sted2576d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2576d,
			Enable=>Enabled2576d,
			match=>matchd2576d,
			run=>run);

	Enabled2576d <= matchd2575d;
	-- d2577d
	sted2577d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2577d,
			Enable=>Enabled2577d,
			match=>matchd2577d,
			run=>run);

	Enabled2577d <= matchd2576d;
	-- d2578d
	sted2578d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2578d,
			Enable=>Enabled2578d,
			match=>matchd2578d,
			run=>run);

	Enabled2578d <= matchd2577d;
	-- d2579d
	sted2579d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2579d,
			Enable=>Enabled2579d,
			match=>matchd2579d,
			run=>run);

	Enabled2579d <= matchd2578d OR matchd2579d;
	-- d2580d
	sted2580d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2580d,
			Enable=>Enabled2580d,
			match=>matchd2580d,
			run=>run);

	Enabled2580d <= matchd2579d;
	-- d2581d
	sted2581d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2581d,
			Enable=>Enabled2581d,
			match=>matchd2581d,
			run=>run);

	Enabled2581d <= matchd2580d;
	-- d2582d
	sted2582d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2582d,
			Enable=>Enabled2582d,
			match=>matchd2582d,
			run=>run);

	Enabled2582d <= matchd2581d;
	-- d2583d
	sted2583d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2583d,
			Enable=>Enabled2583d,
			match=>matchd2583d,
			run=>run);

	Enabled2583d <= matchd2582d;
	-- d2584d
	sted2584d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2584d,
			Enable=>Enabled2584d,
			match=>matchd2584d,
			run=>run);

	Enabled2584d <= matchd2583d OR matchd2584d;
	-- d2585d
	sted2585d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2585d,
			Enable=>Enabled2585d,
			match=>matchd2585d,
			run=>run);

	Enabled2585d <= matchd2584d;
	-- d2586d
	sted2586d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2586d,
			Enable=>Enabled2586d,
			match=>matchd2586d,
			run=>run);

	Enabled2586d <= matchd2585d;
	-- d2587d
	sted2587d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2587d,
			Enable=>Enabled2587d,
			match=>matchd2587d,
			run=>run);

	Enabled2587d <= matchd2586d;
	-- d2588d
	sted2588d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2588d,
			Enable=>Enabled2588d,
			match=>matchd2588d,
			run=>run);

	reports(138) <= matchd2588d;
	Enabled2588d <= matchd2587d;
	-- d2589d
	sted2589d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2589d,
			Enable=>Enabled2589d,
			match=>matchd2589d,
			run=>run);

	-- d2590d
	sted2590d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2590d,
			Enable=>Enabled2590d,
			match=>matchd2590d,
			run=>run);

	Enabled2590d <= matchd2589d OR matchd2590d;
	-- d2591d
	sted2591d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2591d,
			Enable=>Enabled2591d,
			match=>matchd2591d,
			run=>run);

	Enabled2591d <= matchd2590d;
	-- d2592d
	sted2592d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2592d,
			Enable=>Enabled2592d,
			match=>matchd2592d,
			run=>run);

	Enabled2592d <= matchd2591d;
	-- d2593d
	sted2593d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2593d,
			Enable=>Enabled2593d,
			match=>matchd2593d,
			run=>run);

	Enabled2593d <= matchd2592d;
	-- d2594d
	sted2594d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2594d,
			Enable=>Enabled2594d,
			match=>matchd2594d,
			run=>run);

	Enabled2594d <= matchd2593d;
	-- d2595d
	sted2595d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2595d,
			Enable=>Enabled2595d,
			match=>matchd2595d,
			run=>run);

	Enabled2595d <= matchd2594d OR matchd2595d;
	-- d2596d
	sted2596d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2596d,
			Enable=>Enabled2596d,
			match=>matchd2596d,
			run=>run);

	Enabled2596d <= matchd2595d;
	-- d2597d
	sted2597d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2597d,
			Enable=>Enabled2597d,
			match=>matchd2597d,
			run=>run);

	Enabled2597d <= matchd2596d;
	-- d2598d
	sted2598d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2598d,
			Enable=>Enabled2598d,
			match=>matchd2598d,
			run=>run);

	Enabled2598d <= matchd2597d;
	-- d2599d
	sted2599d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2599d,
			Enable=>Enabled2599d,
			match=>matchd2599d,
			run=>run);

	reports(139) <= matchd2599d;
	Enabled2599d <= matchd2598d;
	-- d2600d
	sted2600d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2600d,
			Enable=>Enabled2600d,
			match=>matchd2600d,
			run=>run);

	-- d2601d
	sted2601d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2601d,
			Enable=>Enabled2601d,
			match=>matchd2601d,
			run=>run);

	Enabled2601d <= matchd2600d;
	-- d2602d
	sted2602d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2602d,
			Enable=>Enabled2602d,
			match=>matchd2602d,
			run=>run);

	Enabled2602d <= matchd2601d;
	-- d2603d
	sted2603d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2603d,
			Enable=>Enabled2603d,
			match=>matchd2603d,
			run=>run);

	Enabled2603d <= matchd2602d;
	-- d2604d
	sted2604d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2604d,
			Enable=>Enabled2604d,
			match=>matchd2604d,
			run=>run);

	Enabled2604d <= matchd2603d;
	-- d2605d
	sted2605d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2605d,
			Enable=>Enabled2605d,
			match=>matchd2605d,
			run=>run);

	Enabled2605d <= matchd2604d;
	-- d2606d
	sted2606d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2606d,
			Enable=>Enabled2606d,
			match=>matchd2606d,
			run=>run);

	Enabled2606d <= matchd2605d;
	-- d2607d
	sted2607d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2607d,
			Enable=>Enabled2607d,
			match=>matchd2607d,
			run=>run);

	Enabled2607d <= matchd2606d;
	-- d2608d
	sted2608d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2608d,
			Enable=>Enabled2608d,
			match=>matchd2608d,
			run=>run);

	Enabled2608d <= matchd2607d;
	-- d2609d
	sted2609d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2609d,
			Enable=>Enabled2609d,
			match=>matchd2609d,
			run=>run);

	Enabled2609d <= matchd2608d OR matchd2609d;
	-- d2610d
	sted2610d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2610d,
			Enable=>Enabled2610d,
			match=>matchd2610d,
			run=>run);

	Enabled2610d <= matchd2609d;
	-- d2611d
	sted2611d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2611d,
			Enable=>Enabled2611d,
			match=>matchd2611d,
			run=>run);

	Enabled2611d <= matchd2610d OR matchd2611d;
	-- d2612d
	sted2612d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2612d,
			Enable=>Enabled2612d,
			match=>matchd2612d,
			run=>run);

	Enabled2612d <= matchd2611d;
	-- d2613d
	sted2613d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2613d,
			Enable=>Enabled2613d,
			match=>matchd2613d,
			run=>run);

	Enabled2613d <= matchd2612d OR matchd2613d;
	-- d2614d
	sted2614d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2614d,
			Enable=>Enabled2614d,
			match=>matchd2614d,
			run=>run);

	Enabled2614d <= matchd2613d;
	-- d2615d
	sted2615d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2615d,
			Enable=>Enabled2615d,
			match=>matchd2615d,
			run=>run);

	Enabled2615d <= matchd2614d;
	-- d2616d
	sted2616d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2616d,
			Enable=>Enabled2616d,
			match=>matchd2616d,
			run=>run);

	Enabled2616d <= matchd2615d;
	-- d2617d
	sted2617d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2617d,
			Enable=>Enabled2617d,
			match=>matchd2617d,
			run=>run);

	Enabled2617d <= matchd2616d;
	-- d2618d
	sted2618d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2618d,
			Enable=>Enabled2618d,
			match=>matchd2618d,
			run=>run);

	reports(140) <= matchd2618d;
	Enabled2618d <= matchd2617d;
	-- d2619d
	sted2619d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2619d,
			Enable=>Enabled2619d,
			match=>matchd2619d,
			run=>run);

	-- d2620d
	sted2620d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2620d,
			Enable=>Enabled2620d,
			match=>matchd2620d,
			run=>run);

	Enabled2620d <= matchd2619d OR matchd2620d;
	-- d2621d
	sted2621d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2621d,
			Enable=>Enabled2621d,
			match=>matchd2621d,
			run=>run);

	Enabled2621d <= matchd2620d;
	-- d2622d
	sted2622d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2622d,
			Enable=>Enabled2622d,
			match=>matchd2622d,
			run=>run);

	Enabled2622d <= matchd2621d;
	-- d2623d
	sted2623d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2623d,
			Enable=>Enabled2623d,
			match=>matchd2623d,
			run=>run);

	Enabled2623d <= matchd2622d;
	-- d2624d
	sted2624d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2624d,
			Enable=>Enabled2624d,
			match=>matchd2624d,
			run=>run);

	Enabled2624d <= matchd2623d;
	-- d2625d
	sted2625d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2625d,
			Enable=>Enabled2625d,
			match=>matchd2625d,
			run=>run);

	Enabled2625d <= matchd2624d;
	-- d2626d
	sted2626d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2626d,
			Enable=>Enabled2626d,
			match=>matchd2626d,
			run=>run);

	Enabled2626d <= matchd2626d OR matchd2625d;
	-- d2627d
	sted2627d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2627d,
			Enable=>Enabled2627d,
			match=>matchd2627d,
			run=>run);

	Enabled2627d <= matchd2626d;
	-- d2628d
	sted2628d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2628d,
			Enable=>Enabled2628d,
			match=>matchd2628d,
			run=>run);

	Enabled2628d <= matchd2627d;
	-- d2629d
	sted2629d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2629d,
			Enable=>Enabled2629d,
			match=>matchd2629d,
			run=>run);

	Enabled2629d <= matchd2628d;
	-- d2630d
	sted2630d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2630d,
			Enable=>Enabled2630d,
			match=>matchd2630d,
			run=>run);

	Enabled2630d <= matchd2629d;
	-- d2631d
	sted2631d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2631d,
			Enable=>Enabled2631d,
			match=>matchd2631d,
			run=>run);

	Enabled2631d <= matchd2630d;
	-- d2632d
	sted2632d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2632d,
			Enable=>Enabled2632d,
			match=>matchd2632d,
			run=>run);

	Enabled2632d <= matchd2631d OR matchd2632d;
	-- d2633d
	sted2633d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2633d,
			Enable=>Enabled2633d,
			match=>matchd2633d,
			run=>run);

	Enabled2633d <= matchd2632d;
	-- d2634d
	sted2634d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2634d,
			Enable=>Enabled2634d,
			match=>matchd2634d,
			run=>run);

	Enabled2634d <= matchd2633d;
	-- d2635d
	sted2635d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2635d,
			Enable=>Enabled2635d,
			match=>matchd2635d,
			run=>run);

	reports(141) <= matchd2635d;
	Enabled2635d <= matchd2634d;
	-- d2636d
	sted2636d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2636d,
			Enable=>Enabled2636d,
			match=>matchd2636d,
			run=>run);

	-- d2637d
	sted2637d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2637d,
			Enable=>Enabled2637d,
			match=>matchd2637d,
			run=>run);

	Enabled2637d <= matchd2637d OR matchd2636d;
	-- d2638d
	sted2638d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2638d,
			Enable=>Enabled2638d,
			match=>matchd2638d,
			run=>run);

	Enabled2638d <= matchd2637d;
	-- d2639d
	sted2639d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2639d,
			Enable=>Enabled2639d,
			match=>matchd2639d,
			run=>run);

	Enabled2639d <= matchd2638d;
	-- d2640d
	sted2640d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2640d,
			Enable=>Enabled2640d,
			match=>matchd2640d,
			run=>run);

	Enabled2640d <= matchd2639d;
	-- d2641d
	sted2641d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2641d,
			Enable=>Enabled2641d,
			match=>matchd2641d,
			run=>run);

	Enabled2641d <= matchd2640d;
	-- d2642d
	sted2642d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2642d,
			Enable=>Enabled2642d,
			match=>matchd2642d,
			run=>run);

	Enabled2642d <= matchd2641d OR matchd2642d;
	-- d2643d
	sted2643d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2643d,
			Enable=>Enabled2643d,
			match=>matchd2643d,
			run=>run);

	Enabled2643d <= matchd2642d;
	-- d2644d
	sted2644d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2644d,
			Enable=>Enabled2644d,
			match=>matchd2644d,
			run=>run);

	Enabled2644d <= matchd2643d;
	-- d2645d
	sted2645d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2645d,
			Enable=>Enabled2645d,
			match=>matchd2645d,
			run=>run);

	Enabled2645d <= matchd2644d;
	-- d2646d
	sted2646d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2646d,
			Enable=>Enabled2646d,
			match=>matchd2646d,
			run=>run);

	Enabled2646d <= matchd2645d;
	-- d2647d
	sted2647d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2647d,
			Enable=>Enabled2647d,
			match=>matchd2647d,
			run=>run);

	reports(142) <= matchd2647d;
	Enabled2647d <= matchd2646d;
	-- d2648d
	sted2648d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2648d,
			Enable=>Enabled2648d,
			match=>matchd2648d,
			run=>run);

	-- d2649d
	sted2649d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2649d,
			Enable=>Enabled2649d,
			match=>matchd2649d,
			run=>run);

	Enabled2649d <= matchd2648d OR matchd2649d;
	-- d2650d
	sted2650d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2650d,
			Enable=>Enabled2650d,
			match=>matchd2650d,
			run=>run);

	Enabled2650d <= matchd2649d;
	-- d2651d
	sted2651d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2651d,
			Enable=>Enabled2651d,
			match=>matchd2651d,
			run=>run);

	Enabled2651d <= matchd2650d;
	-- d2652d
	sted2652d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2652d,
			Enable=>Enabled2652d,
			match=>matchd2652d,
			run=>run);

	Enabled2652d <= matchd2651d;
	-- d2653d
	sted2653d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2653d,
			Enable=>Enabled2653d,
			match=>matchd2653d,
			run=>run);

	Enabled2653d <= matchd2652d;
	-- d2654d
	sted2654d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2654d,
			Enable=>Enabled2654d,
			match=>matchd2654d,
			run=>run);

	Enabled2654d <= matchd2654d OR matchd2653d;
	-- d2655d
	sted2655d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2655d,
			Enable=>Enabled2655d,
			match=>matchd2655d,
			run=>run);

	Enabled2655d <= matchd2654d;
	-- d2656d
	sted2656d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2656d,
			Enable=>Enabled2656d,
			match=>matchd2656d,
			run=>run);

	Enabled2656d <= matchd2655d;
	-- d2657d
	sted2657d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2657d,
			Enable=>Enabled2657d,
			match=>matchd2657d,
			run=>run);

	Enabled2657d <= matchd2656d;
	-- d2658d
	sted2658d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2658d,
			Enable=>Enabled2658d,
			match=>matchd2658d,
			run=>run);

	Enabled2658d <= matchd2657d;
	-- d2659d
	sted2659d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2659d,
			Enable=>Enabled2659d,
			match=>matchd2659d,
			run=>run);

	reports(143) <= matchd2659d;
	Enabled2659d <= matchd2658d;
	-- d2660d
	sted2660d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2660d,
			Enable=>Enabled2660d,
			match=>matchd2660d,
			run=>run);

	-- d2661d
	sted2661d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2661d,
			Enable=>Enabled2661d,
			match=>matchd2661d,
			run=>run);

	Enabled2661d <= matchd2660d OR matchd2661d;
	-- d2662d
	sted2662d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2662d,
			Enable=>Enabled2662d,
			match=>matchd2662d,
			run=>run);

	Enabled2662d <= matchd2661d;
	-- d2663d
	sted2663d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2663d,
			Enable=>Enabled2663d,
			match=>matchd2663d,
			run=>run);

	Enabled2663d <= matchd2662d;
	-- d2664d
	sted2664d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2664d,
			Enable=>Enabled2664d,
			match=>matchd2664d,
			run=>run);

	Enabled2664d <= matchd2663d;
	-- d2665d
	sted2665d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2665d,
			Enable=>Enabled2665d,
			match=>matchd2665d,
			run=>run);

	Enabled2665d <= matchd2664d;
	-- d2666d
	sted2666d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2666d,
			Enable=>Enabled2666d,
			match=>matchd2666d,
			run=>run);

	Enabled2666d <= matchd2666d OR matchd2665d;
	-- d2667d
	sted2667d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2667d,
			Enable=>Enabled2667d,
			match=>matchd2667d,
			run=>run);

	Enabled2667d <= matchd2666d;
	-- d2668d
	sted2668d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2668d,
			Enable=>Enabled2668d,
			match=>matchd2668d,
			run=>run);

	Enabled2668d <= matchd2667d;
	-- d2669d
	sted2669d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2669d,
			Enable=>Enabled2669d,
			match=>matchd2669d,
			run=>run);

	Enabled2669d <= matchd2668d;
	-- d2670d
	sted2670d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2670d,
			Enable=>Enabled2670d,
			match=>matchd2670d,
			run=>run);

	Enabled2670d <= matchd2669d;
	-- d2671d
	sted2671d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2671d,
			Enable=>Enabled2671d,
			match=>matchd2671d,
			run=>run);

	reports(144) <= matchd2671d;
	Enabled2671d <= matchd2670d;
	-- d2672d
	sted2672d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2672d,
			Enable=>Enabled2672d,
			match=>matchd2672d,
			run=>run);

	-- d2673d
	sted2673d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2673d,
			Enable=>Enabled2673d,
			match=>matchd2673d,
			run=>run);

	Enabled2673d <= matchd2673d OR matchd2672d;
	-- d2674d
	sted2674d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2674d,
			Enable=>Enabled2674d,
			match=>matchd2674d,
			run=>run);

	Enabled2674d <= matchd2673d;
	-- d2675d
	sted2675d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2675d,
			Enable=>Enabled2675d,
			match=>matchd2675d,
			run=>run);

	Enabled2675d <= matchd2674d;
	-- d2676d
	sted2676d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2676d,
			Enable=>Enabled2676d,
			match=>matchd2676d,
			run=>run);

	Enabled2676d <= matchd2675d;
	-- d2677d
	sted2677d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2677d,
			Enable=>Enabled2677d,
			match=>matchd2677d,
			run=>run);

	Enabled2677d <= matchd2676d;
	-- d2678d
	sted2678d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2678d,
			Enable=>Enabled2678d,
			match=>matchd2678d,
			run=>run);

	Enabled2678d <= matchd2677d OR matchd2678d;
	-- d2679d
	sted2679d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2679d,
			Enable=>Enabled2679d,
			match=>matchd2679d,
			run=>run);

	Enabled2679d <= matchd2678d;
	-- d2680d
	sted2680d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2680d,
			Enable=>Enabled2680d,
			match=>matchd2680d,
			run=>run);

	Enabled2680d <= matchd2679d;
	-- d2681d
	sted2681d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2681d,
			Enable=>Enabled2681d,
			match=>matchd2681d,
			run=>run);

	Enabled2681d <= matchd2680d;
	-- d2682d
	sted2682d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2682d,
			Enable=>Enabled2682d,
			match=>matchd2682d,
			run=>run);

	Enabled2682d <= matchd2681d;
	-- d2683d
	sted2683d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2683d,
			Enable=>Enabled2683d,
			match=>matchd2683d,
			run=>run);

	Enabled2683d <= matchd2682d OR matchd2683d;
	-- d2684d
	sted2684d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2684d,
			Enable=>Enabled2684d,
			match=>matchd2684d,
			run=>run);

	Enabled2684d <= matchd2683d;
	-- d2685d
	sted2685d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2685d,
			Enable=>Enabled2685d,
			match=>matchd2685d,
			run=>run);

	Enabled2685d <= matchd2684d;
	-- d2686d
	sted2686d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2686d,
			Enable=>Enabled2686d,
			match=>matchd2686d,
			run=>run);

	Enabled2686d <= matchd2685d;
	-- d2687d
	sted2687d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2687d,
			Enable=>Enabled2687d,
			match=>matchd2687d,
			run=>run);

	reports(145) <= matchd2687d;
	Enabled2687d <= matchd2686d;
	-- d2688d
	sted2688d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2688d,
			Enable=>Enabled2688d,
			match=>matchd2688d,
			run=>run);

	-- d2689d
	sted2689d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2689d,
			Enable=>Enabled2689d,
			match=>matchd2689d,
			run=>run);

	Enabled2689d <= matchd2688d;
	-- d2690d
	sted2690d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2690d,
			Enable=>Enabled2690d,
			match=>matchd2690d,
			run=>run);

	Enabled2690d <= matchd2689d;
	-- d2691d
	sted2691d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2691d,
			Enable=>Enabled2691d,
			match=>matchd2691d,
			run=>run);

	Enabled2691d <= matchd2690d;
	-- d2692d
	sted2692d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2692d,
			Enable=>Enabled2692d,
			match=>matchd2692d,
			run=>run);

	Enabled2692d <= matchd2691d;
	-- d2693d
	sted2693d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2693d,
			Enable=>Enabled2693d,
			match=>matchd2693d,
			run=>run);

	Enabled2693d <= matchd2692d;
	-- d2694d
	sted2694d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2694d,
			Enable=>Enabled2694d,
			match=>matchd2694d,
			run=>run);

	Enabled2694d <= matchd2693d;
	-- d2695d
	sted2695d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2695d,
			Enable=>Enabled2695d,
			match=>matchd2695d,
			run=>run);

	Enabled2695d <= matchd2694d;
	-- d2696d
	sted2696d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2696d,
			Enable=>Enabled2696d,
			match=>matchd2696d,
			run=>run);

	Enabled2696d <= matchd2695d;
	-- d2697d
	sted2697d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2697d,
			Enable=>Enabled2697d,
			match=>matchd2697d,
			run=>run);

	reports(146) <= matchd2697d;
	Enabled2697d <= matchd2696d;
	-- d2698d
	sted2698d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2698d,
			Enable=>Enabled2698d,
			match=>matchd2698d,
			run=>run);

	-- d2699d
	sted2699d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2699d,
			Enable=>Enabled2699d,
			match=>matchd2699d,
			run=>run);

	Enabled2699d <= matchd2699d OR matchd2698d;
	-- d2700d
	sted2700d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2700d,
			Enable=>Enabled2700d,
			match=>matchd2700d,
			run=>run);

	Enabled2700d <= matchd2699d;
	-- d2701d
	sted2701d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2701d,
			Enable=>Enabled2701d,
			match=>matchd2701d,
			run=>run);

	Enabled2701d <= matchd2700d;
	-- d2702d
	sted2702d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2702d,
			Enable=>Enabled2702d,
			match=>matchd2702d,
			run=>run);

	Enabled2702d <= matchd2701d;
	-- d2703d
	sted2703d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2703d,
			Enable=>Enabled2703d,
			match=>matchd2703d,
			run=>run);

	Enabled2703d <= matchd2702d;
	-- d2704d
	sted2704d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2704d,
			Enable=>Enabled2704d,
			match=>matchd2704d,
			run=>run);

	Enabled2704d <= matchd2703d OR matchd2704d;
	-- d2705d
	sted2705d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2705d,
			Enable=>Enabled2705d,
			match=>matchd2705d,
			run=>run);

	Enabled2705d <= matchd2704d;
	-- d2706d
	sted2706d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2706d,
			Enable=>Enabled2706d,
			match=>matchd2706d,
			run=>run);

	Enabled2706d <= matchd2705d;
	-- d2707d
	sted2707d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2707d,
			Enable=>Enabled2707d,
			match=>matchd2707d,
			run=>run);

	Enabled2707d <= matchd2706d;
	-- d2708d
	sted2708d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2708d,
			Enable=>Enabled2708d,
			match=>matchd2708d,
			run=>run);

	Enabled2708d <= matchd2707d;
	-- d2709d
	sted2709d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2709d,
			Enable=>Enabled2709d,
			match=>matchd2709d,
			run=>run);

	Enabled2709d <= matchd2709d OR matchd2708d;
	-- d2710d
	sted2710d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2710d,
			Enable=>Enabled2710d,
			match=>matchd2710d,
			run=>run);

	Enabled2710d <= matchd2709d;
	-- d2711d
	sted2711d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2711d,
			Enable=>Enabled2711d,
			match=>matchd2711d,
			run=>run);

	Enabled2711d <= matchd2710d;
	-- d2712d
	sted2712d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2712d,
			Enable=>Enabled2712d,
			match=>matchd2712d,
			run=>run);

	reports(147) <= matchd2712d;
	Enabled2712d <= matchd2711d;
	-- d2713d
	sted2713d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2713d,
			Enable=>Enabled2713d,
			match=>matchd2713d,
			run=>run);

	-- d2714d
	sted2714d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2714d,
			Enable=>Enabled2714d,
			match=>matchd2714d,
			run=>run);

	Enabled2714d <= matchd2713d;
	-- d2715d
	sted2715d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2715d,
			Enable=>Enabled2715d,
			match=>matchd2715d,
			run=>run);

	Enabled2715d <= matchd2714d;
	-- d2716d
	sted2716d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2716d,
			Enable=>Enabled2716d,
			match=>matchd2716d,
			run=>run);

	Enabled2716d <= matchd2715d;
	-- d2717d
	sted2717d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2717d,
			Enable=>Enabled2717d,
			match=>matchd2717d,
			run=>run);

	Enabled2717d <= matchd2716d;
	-- d2718d
	sted2718d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2718d,
			Enable=>Enabled2718d,
			match=>matchd2718d,
			run=>run);

	Enabled2718d <= matchd2717d;
	-- d2719d
	sted2719d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2719d,
			Enable=>Enabled2719d,
			match=>matchd2719d,
			run=>run);

	Enabled2719d <= matchd2718d;
	-- d2720d
	sted2720d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2720d,
			Enable=>Enabled2720d,
			match=>matchd2720d,
			run=>run);

	reports(148) <= matchd2720d;
	Enabled2720d <= matchd2719d;
	-- d2721d
	sted2721d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2721d,
			Enable=>Enabled2721d,
			match=>matchd2721d,
			run=>run);

	-- d2722d
	sted2722d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2722d,
			Enable=>Enabled2722d,
			match=>matchd2722d,
			run=>run);

	Enabled2722d <= matchd2722d OR matchd2721d;
	-- d2723d
	sted2723d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2723d,
			Enable=>Enabled2723d,
			match=>matchd2723d,
			run=>run);

	Enabled2723d <= matchd2722d;
	-- d2724d
	sted2724d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2724d,
			Enable=>Enabled2724d,
			match=>matchd2724d,
			run=>run);

	Enabled2724d <= matchd2723d;
	-- d2725d
	sted2725d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2725d,
			Enable=>Enabled2725d,
			match=>matchd2725d,
			run=>run);

	Enabled2725d <= matchd2724d;
	-- d2726d
	sted2726d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2726d,
			Enable=>Enabled2726d,
			match=>matchd2726d,
			run=>run);

	Enabled2726d <= matchd2725d;
	-- d2727d
	sted2727d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2727d,
			Enable=>Enabled2727d,
			match=>matchd2727d,
			run=>run);

	Enabled2727d <= matchd2726d;
	-- d2728d
	sted2728d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2728d,
			Enable=>Enabled2728d,
			match=>matchd2728d,
			run=>run);

	Enabled2728d <= matchd2727d;
	-- d2729d
	sted2729d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2729d,
			Enable=>Enabled2729d,
			match=>matchd2729d,
			run=>run);

	Enabled2729d <= matchd2728d;
	-- d2730d
	sted2730d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2730d,
			Enable=>Enabled2730d,
			match=>matchd2730d,
			run=>run);

	Enabled2730d <= matchd2729d;
	-- d2731d
	sted2731d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2731d,
			Enable=>Enabled2731d,
			match=>matchd2731d,
			run=>run);

	Enabled2731d <= matchd2730d OR matchd2731d;
	-- d2732d
	sted2732d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2732d,
			Enable=>Enabled2732d,
			match=>matchd2732d,
			run=>run);

	Enabled2732d <= matchd2731d;
	-- d2733d
	sted2733d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2733d,
			Enable=>Enabled2733d,
			match=>matchd2733d,
			run=>run);

	Enabled2733d <= matchd2732d;
	-- d2734d
	sted2734d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2734d,
			Enable=>Enabled2734d,
			match=>matchd2734d,
			run=>run);

	Enabled2734d <= matchd2733d;
	-- d2735d
	sted2735d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2735d,
			Enable=>Enabled2735d,
			match=>matchd2735d,
			run=>run);

	Enabled2735d <= matchd2734d;
	-- d2736d
	sted2736d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2736d,
			Enable=>Enabled2736d,
			match=>matchd2736d,
			run=>run);

	Enabled2736d <= matchd2735d;
	-- d2737d
	sted2737d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2737d,
			Enable=>Enabled2737d,
			match=>matchd2737d,
			run=>run);

	Enabled2737d <= matchd2736d OR matchd2737d;
	-- d2738d
	sted2738d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2738d,
			Enable=>Enabled2738d,
			match=>matchd2738d,
			run=>run);

	Enabled2738d <= matchd2737d;
	-- d2739d
	sted2739d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2739d,
			Enable=>Enabled2739d,
			match=>matchd2739d,
			run=>run);

	Enabled2739d <= matchd2738d;
	-- d2740d
	sted2740d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2740d,
			Enable=>Enabled2740d,
			match=>matchd2740d,
			run=>run);

	Enabled2740d <= matchd2739d;
	-- d2741d
	sted2741d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2741d,
			Enable=>Enabled2741d,
			match=>matchd2741d,
			run=>run);

	reports(149) <= matchd2741d;
	Enabled2741d <= matchd2740d;
	-- d2742d
	sted2742d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2742d,
			Enable=>Enabled2742d,
			match=>matchd2742d,
			run=>run);

	-- d2743d
	sted2743d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2743d,
			Enable=>Enabled2743d,
			match=>matchd2743d,
			run=>run);

	Enabled2743d <= matchd2742d OR matchd2743d;
	-- d2744d
	sted2744d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2744d,
			Enable=>Enabled2744d,
			match=>matchd2744d,
			run=>run);

	Enabled2744d <= matchd2743d;
	-- d2745d
	sted2745d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2745d,
			Enable=>Enabled2745d,
			match=>matchd2745d,
			run=>run);

	Enabled2745d <= matchd2744d;
	-- d2746d
	sted2746d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2746d,
			Enable=>Enabled2746d,
			match=>matchd2746d,
			run=>run);

	Enabled2746d <= matchd2745d;
	-- d2747d
	sted2747d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2747d,
			Enable=>Enabled2747d,
			match=>matchd2747d,
			run=>run);

	Enabled2747d <= matchd2746d;
	-- d2748d
	sted2748d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2748d,
			Enable=>Enabled2748d,
			match=>matchd2748d,
			run=>run);

	Enabled2748d <= matchd2747d;
	-- d2749d
	sted2749d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2749d,
			Enable=>Enabled2749d,
			match=>matchd2749d,
			run=>run);

	Enabled2749d <= matchd2748d;
	-- d2750d
	sted2750d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2750d,
			Enable=>Enabled2750d,
			match=>matchd2750d,
			run=>run);

	Enabled2750d <= matchd2749d;
	-- d2751d
	sted2751d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2751d,
			Enable=>Enabled2751d,
			match=>matchd2751d,
			run=>run);

	Enabled2751d <= matchd2750d;
	-- d2752d
	sted2752d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2752d,
			Enable=>Enabled2752d,
			match=>matchd2752d,
			run=>run);

	Enabled2752d <= matchd2751d OR matchd2752d;
	-- d2753d
	sted2753d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2753d,
			Enable=>Enabled2753d,
			match=>matchd2753d,
			run=>run);

	Enabled2753d <= matchd2752d;
	-- d2754d
	sted2754d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2754d,
			Enable=>Enabled2754d,
			match=>matchd2754d,
			run=>run);

	Enabled2754d <= matchd2753d;
	-- d2755d
	sted2755d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2755d,
			Enable=>Enabled2755d,
			match=>matchd2755d,
			run=>run);

	Enabled2755d <= matchd2754d;
	-- d2756d
	sted2756d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2756d,
			Enable=>Enabled2756d,
			match=>matchd2756d,
			run=>run);

	Enabled2756d <= matchd2755d;
	-- d2757d
	sted2757d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2757d,
			Enable=>Enabled2757d,
			match=>matchd2757d,
			run=>run);

	Enabled2757d <= matchd2756d;
	-- d2758d
	sted2758d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2758d,
			Enable=>Enabled2758d,
			match=>matchd2758d,
			run=>run);

	Enabled2758d <= matchd2757d OR matchd2758d;
	-- d2759d
	sted2759d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2759d,
			Enable=>Enabled2759d,
			match=>matchd2759d,
			run=>run);

	Enabled2759d <= matchd2758d;
	-- d2760d
	sted2760d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2760d,
			Enable=>Enabled2760d,
			match=>matchd2760d,
			run=>run);

	Enabled2760d <= matchd2759d;
	-- d2761d
	sted2761d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2761d,
			Enable=>Enabled2761d,
			match=>matchd2761d,
			run=>run);

	Enabled2761d <= matchd2760d;
	-- d2762d
	sted2762d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2762d,
			Enable=>Enabled2762d,
			match=>matchd2762d,
			run=>run);

	reports(150) <= matchd2762d;
	Enabled2762d <= matchd2761d;
	-- d2763d
	sted2763d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2763d,
			Enable=>Enabled2763d,
			match=>matchd2763d,
			run=>run);

	-- d2764d
	sted2764d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2764d,
			Enable=>Enabled2764d,
			match=>matchd2764d,
			run=>run);

	Enabled2764d <= matchd2763d;
	-- d2765d
	sted2765d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2765d,
			Enable=>Enabled2765d,
			match=>matchd2765d,
			run=>run);

	Enabled2765d <= matchd2764d;
	-- d2766d
	sted2766d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2766d,
			Enable=>Enabled2766d,
			match=>matchd2766d,
			run=>run);

	Enabled2766d <= matchd2765d;
	-- d2767d
	sted2767d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2767d,
			Enable=>Enabled2767d,
			match=>matchd2767d,
			run=>run);

	Enabled2767d <= matchd2766d;
	-- d2768d
	sted2768d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2768d,
			Enable=>Enabled2768d,
			match=>matchd2768d,
			run=>run);

	Enabled2768d <= matchd2767d;
	-- d2769d
	sted2769d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2769d,
			Enable=>Enabled2769d,
			match=>matchd2769d,
			run=>run);

	Enabled2769d <= matchd2768d;
	-- d2770d
	sted2770d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2770d,
			Enable=>Enabled2770d,
			match=>matchd2770d,
			run=>run);

	Enabled2770d <= matchd2769d;
	-- d2771d
	sted2771d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2771d,
			Enable=>Enabled2771d,
			match=>matchd2771d,
			run=>run);

	Enabled2771d <= matchd2770d;
	-- d2772d
	sted2772d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2772d,
			Enable=>Enabled2772d,
			match=>matchd2772d,
			run=>run);

	Enabled2772d <= matchd2771d;
	-- d2773d
	sted2773d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2773d,
			Enable=>Enabled2773d,
			match=>matchd2773d,
			run=>run);

	Enabled2773d <= matchd2772d;
	-- d2774d
	sted2774d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2774d,
			Enable=>Enabled2774d,
			match=>matchd2774d,
			run=>run);

	Enabled2774d <= matchd2773d;
	-- d2775d
	sted2775d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2775d,
			Enable=>Enabled2775d,
			match=>matchd2775d,
			run=>run);

	reports(151) <= matchd2775d;
	Enabled2775d <= matchd2774d;
	-- d2776d
	sted2776d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2776d,
			Enable=>Enabled2776d,
			match=>matchd2776d,
			run=>run);

	-- d2777d
	sted2777d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2777d,
			Enable=>Enabled2777d,
			match=>matchd2777d,
			run=>run);

	Enabled2777d <= matchd2776d;
	-- d2778d
	sted2778d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2778d,
			Enable=>Enabled2778d,
			match=>matchd2778d,
			run=>run);

	Enabled2778d <= matchd2777d;
	-- d2779d
	sted2779d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2779d,
			Enable=>Enabled2779d,
			match=>matchd2779d,
			run=>run);

	Enabled2779d <= matchd2778d;
	-- d2780d
	sted2780d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2780d,
			Enable=>Enabled2780d,
			match=>matchd2780d,
			run=>run);

	Enabled2780d <= matchd2779d;
	-- d2781d
	sted2781d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2781d,
			Enable=>Enabled2781d,
			match=>matchd2781d,
			run=>run);

	Enabled2781d <= matchd2780d;
	-- d2782d
	sted2782d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2782d,
			Enable=>Enabled2782d,
			match=>matchd2782d,
			run=>run);

	Enabled2782d <= matchd2781d;
	-- d2783d
	sted2783d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2783d,
			Enable=>Enabled2783d,
			match=>matchd2783d,
			run=>run);

	Enabled2783d <= matchd2782d;
	-- d2784d
	sted2784d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2784d,
			Enable=>Enabled2784d,
			match=>matchd2784d,
			run=>run);

	Enabled2784d <= matchd2783d;
	-- d2785d
	sted2785d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2785d,
			Enable=>Enabled2785d,
			match=>matchd2785d,
			run=>run);

	Enabled2785d <= matchd2784d;
	-- d2786d
	sted2786d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2786d,
			Enable=>Enabled2786d,
			match=>matchd2786d,
			run=>run);

	Enabled2786d <= matchd2786d OR matchd2785d;
	-- d2787d
	sted2787d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2787d,
			Enable=>Enabled2787d,
			match=>matchd2787d,
			run=>run);

	Enabled2787d <= matchd2786d;
	-- d2788d
	sted2788d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2788d,
			Enable=>Enabled2788d,
			match=>matchd2788d,
			run=>run);

	Enabled2788d <= matchd2787d;
	-- d2789d
	sted2789d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2789d,
			Enable=>Enabled2789d,
			match=>matchd2789d,
			run=>run);

	Enabled2789d <= matchd2788d;
	-- d2790d
	sted2790d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2790d,
			Enable=>Enabled2790d,
			match=>matchd2790d,
			run=>run);

	reports(152) <= matchd2790d;
	Enabled2790d <= matchd2789d;
	-- d2791d
	sted2791d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2791d,
			Enable=>Enabled2791d,
			match=>matchd2791d,
			run=>run);

	-- d2792d
	sted2792d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2792d,
			Enable=>Enabled2792d,
			match=>matchd2792d,
			run=>run);

	Enabled2792d <= matchd2792d OR matchd2791d;
	-- d2793d
	sted2793d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2793d,
			Enable=>Enabled2793d,
			match=>matchd2793d,
			run=>run);

	Enabled2793d <= matchd2792d;
	-- d2794d
	sted2794d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2794d,
			Enable=>Enabled2794d,
			match=>matchd2794d,
			run=>run);

	Enabled2794d <= matchd2793d;
	-- d2795d
	sted2795d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2795d,
			Enable=>Enabled2795d,
			match=>matchd2795d,
			run=>run);

	Enabled2795d <= matchd2794d;
	-- d2796d
	sted2796d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2796d,
			Enable=>Enabled2796d,
			match=>matchd2796d,
			run=>run);

	Enabled2796d <= matchd2795d;
	-- d2797d
	sted2797d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2797d,
			Enable=>Enabled2797d,
			match=>matchd2797d,
			run=>run);

	Enabled2797d <= matchd2796d OR matchd2797d;
	-- d2798d
	sted2798d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2798d,
			Enable=>Enabled2798d,
			match=>matchd2798d,
			run=>run);

	Enabled2798d <= matchd2797d;
	-- d2799d
	sted2799d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2799d,
			Enable=>Enabled2799d,
			match=>matchd2799d,
			run=>run);

	Enabled2799d <= matchd2798d;
	-- d2800d
	sted2800d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2800d,
			Enable=>Enabled2800d,
			match=>matchd2800d,
			run=>run);

	Enabled2800d <= matchd2799d;
	-- d2801d
	sted2801d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2801d,
			Enable=>Enabled2801d,
			match=>matchd2801d,
			run=>run);

	reports(153) <= matchd2801d;
	Enabled2801d <= matchd2800d;
	-- d2802d
	sted2802d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2802d,
			Enable=>Enabled2802d,
			match=>matchd2802d,
			run=>run);

	-- d2803d
	sted2803d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2803d,
			Enable=>Enabled2803d,
			match=>matchd2803d,
			run=>run);

	Enabled2803d <= matchd2803d OR matchd2802d;
	-- d2804d
	sted2804d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2804d,
			Enable=>Enabled2804d,
			match=>matchd2804d,
			run=>run);

	Enabled2804d <= matchd2803d;
	-- d2805d
	sted2805d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2805d,
			Enable=>Enabled2805d,
			match=>matchd2805d,
			run=>run);

	Enabled2805d <= matchd2804d OR matchd2805d;
	-- d2806d
	sted2806d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2806d,
			Enable=>Enabled2806d,
			match=>matchd2806d,
			run=>run);

	Enabled2806d <= matchd2805d;
	-- d2807d
	sted2807d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2807d,
			Enable=>Enabled2807d,
			match=>matchd2807d,
			run=>run);

	Enabled2807d <= matchd2806d OR matchd2807d;
	-- d2808d
	sted2808d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2808d,
			Enable=>Enabled2808d,
			match=>matchd2808d,
			run=>run);

	Enabled2808d <= matchd2807d;
	-- d2809d
	sted2809d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2809d,
			Enable=>Enabled2809d,
			match=>matchd2809d,
			run=>run);

	Enabled2809d <= matchd2808d;
	-- d2810d
	sted2810d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2810d,
			Enable=>Enabled2810d,
			match=>matchd2810d,
			run=>run);

	Enabled2810d <= matchd2809d;
	-- d2811d
	sted2811d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2811d,
			Enable=>Enabled2811d,
			match=>matchd2811d,
			run=>run);

	Enabled2811d <= matchd2810d;
	-- d2812d
	sted2812d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2812d,
			Enable=>Enabled2812d,
			match=>matchd2812d,
			run=>run);

	Enabled2812d <= matchd2811d;
	-- d2813d
	sted2813d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2813d,
			Enable=>Enabled2813d,
			match=>matchd2813d,
			run=>run);

	Enabled2813d <= matchd2813d OR matchd2812d;
	-- d2814d
	sted2814d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2814d,
			Enable=>Enabled2814d,
			match=>matchd2814d,
			run=>run);

	Enabled2814d <= matchd2813d;
	-- d2815d
	sted2815d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2815d,
			Enable=>Enabled2815d,
			match=>matchd2815d,
			run=>run);

	Enabled2815d <= matchd2814d;
	-- d2816d
	sted2816d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2816d,
			Enable=>Enabled2816d,
			match=>matchd2816d,
			run=>run);

	Enabled2816d <= matchd2815d;
	-- d2817d
	sted2817d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2817d,
			Enable=>Enabled2817d,
			match=>matchd2817d,
			run=>run);

	Enabled2817d <= matchd2816d;
	-- d2818d
	sted2818d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2818d,
			Enable=>Enabled2818d,
			match=>matchd2818d,
			run=>run);

	Enabled2818d <= matchd2817d;
	-- d2819d
	sted2819d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2819d,
			Enable=>Enabled2819d,
			match=>matchd2819d,
			run=>run);

	-- d2820d
	sted2820d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2820d,
			Enable=>Enabled2820d,
			match=>matchd2820d,
			run=>run);

	Enabled2820d <= matchd2820d OR matchd2819d;
	-- d2821d
	sted2821d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2821d,
			Enable=>Enabled2821d,
			match=>matchd2821d,
			run=>run);

	Enabled2821d <= matchd2820d;
	-- d2822d
	sted2822d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2822d,
			Enable=>Enabled2822d,
			match=>matchd2822d,
			run=>run);

	Enabled2822d <= matchd2821d;
	-- d2823d
	sted2823d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2823d,
			Enable=>Enabled2823d,
			match=>matchd2823d,
			run=>run);

	Enabled2823d <= matchd2822d;
	-- d2824d
	sted2824d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2824d,
			Enable=>Enabled2824d,
			match=>matchd2824d,
			run=>run);

	Enabled2824d <= matchd2823d;
	-- d2825d
	sted2825d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2825d,
			Enable=>Enabled2825d,
			match=>matchd2825d,
			run=>run);

	Enabled2825d <= matchd2824d;
	-- d2826d
	sted2826d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2826d,
			Enable=>Enabled2826d,
			match=>matchd2826d,
			run=>run);

	Enabled2826d <= matchd2826d OR matchd2825d;
	-- d2827d
	sted2827d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2827d,
			Enable=>Enabled2827d,
			match=>matchd2827d,
			run=>run);

	Enabled2827d <= matchd2826d;
	-- d2828d
	sted2828d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2828d,
			Enable=>Enabled2828d,
			match=>matchd2828d,
			run=>run);

	Enabled2828d <= matchd2827d OR matchd2828d;
	-- d2829d
	sted2829d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2829d,
			Enable=>Enabled2829d,
			match=>matchd2829d,
			run=>run);

	Enabled2829d <= matchd2828d;
	-- d2830d
	sted2830d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2830d,
			Enable=>Enabled2830d,
			match=>matchd2830d,
			run=>run);

	Enabled2830d <= matchd2830d OR matchd2829d;
	-- d2831d
	sted2831d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2831d,
			Enable=>Enabled2831d,
			match=>matchd2831d,
			run=>run);

	Enabled2831d <= matchd2830d;
	-- d2832d
	sted2832d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2832d,
			Enable=>Enabled2832d,
			match=>matchd2832d,
			run=>run);

	Enabled2832d <= matchd2831d;
	-- d2833d
	sted2833d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2833d,
			Enable=>Enabled2833d,
			match=>matchd2833d,
			run=>run);

	Enabled2833d <= matchd2832d;
	-- d2834d
	sted2834d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2834d,
			Enable=>Enabled2834d,
			match=>matchd2834d,
			run=>run);

	Enabled2834d <= matchd2833d;
	-- d2835d
	sted2835d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2835d,
			Enable=>Enabled2835d,
			match=>matchd2835d,
			run=>run);

	Enabled2835d <= matchd2834d;
	-- d2837d
	sted2837d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2837d,
			Enable=>Enabled2837d,
			match=>matchd2837d,
			run=>run);

	-- d2838d
	sted2838d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2838d,
			Enable=>Enabled2838d,
			match=>matchd2838d,
			run=>run);

	Enabled2838d <= matchd2838d OR matchd2837d;
	-- d2839d
	sted2839d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2839d,
			Enable=>Enabled2839d,
			match=>matchd2839d,
			run=>run);

	Enabled2839d <= matchd2838d;
	-- d2840d
	sted2840d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2840d,
			Enable=>Enabled2840d,
			match=>matchd2840d,
			run=>run);

	Enabled2840d <= matchd2839d;
	-- d2841d
	sted2841d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2841d,
			Enable=>Enabled2841d,
			match=>matchd2841d,
			run=>run);

	Enabled2841d <= matchd2840d;
	-- d2842d
	sted2842d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2842d,
			Enable=>Enabled2842d,
			match=>matchd2842d,
			run=>run);

	Enabled2842d <= matchd2841d;
	-- d2843d
	sted2843d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2843d,
			Enable=>Enabled2843d,
			match=>matchd2843d,
			run=>run);

	Enabled2843d <= matchd2843d OR matchd2842d;
	-- d2844d
	sted2844d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2844d,
			Enable=>Enabled2844d,
			match=>matchd2844d,
			run=>run);

	Enabled2844d <= matchd2843d;
	-- d2845d
	sted2845d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2845d,
			Enable=>Enabled2845d,
			match=>matchd2845d,
			run=>run);

	Enabled2845d <= matchd2844d;
	-- d2846d
	sted2846d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2846d,
			Enable=>Enabled2846d,
			match=>matchd2846d,
			run=>run);

	Enabled2846d <= matchd2845d;
	-- d2847d
	sted2847d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2847d,
			Enable=>Enabled2847d,
			match=>matchd2847d,
			run=>run);

	Enabled2847d <= matchd2846d;
	-- d2848d
	sted2848d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2848d,
			Enable=>Enabled2848d,
			match=>matchd2848d,
			run=>run);

	Enabled2848d <= matchd2847d;
	-- d2849d
	sted2849d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2849d,
			Enable=>Enabled2849d,
			match=>matchd2849d,
			run=>run);

	Enabled2849d <= matchd2849d OR matchd2848d;
	-- d2850d
	sted2850d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2850d,
			Enable=>Enabled2850d,
			match=>matchd2850d,
			run=>run);

	Enabled2850d <= matchd2849d;
	-- d2851d
	sted2851d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2851d,
			Enable=>Enabled2851d,
			match=>matchd2851d,
			run=>run);

	Enabled2851d <= matchd2850d OR matchd2851d;
	-- d2852d
	sted2852d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2852d,
			Enable=>Enabled2852d,
			match=>matchd2852d,
			run=>run);

	Enabled2852d <= matchd2851d;
	-- d2853d
	sted2853d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2853d,
			Enable=>Enabled2853d,
			match=>matchd2853d,
			run=>run);

	-- d2854d
	sted2854d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2854d,
			Enable=>Enabled2854d,
			match=>matchd2854d,
			run=>run);

	Enabled2854d <= matchd2853d OR matchd2854d;
	-- d2855d
	sted2855d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2855d,
			Enable=>Enabled2855d,
			match=>matchd2855d,
			run=>run);

	Enabled2855d <= matchd2854d;
	-- d2856d
	sted2856d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2856d,
			Enable=>Enabled2856d,
			match=>matchd2856d,
			run=>run);

	Enabled2856d <= matchd2855d;
	-- d2857d
	sted2857d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2857d,
			Enable=>Enabled2857d,
			match=>matchd2857d,
			run=>run);

	Enabled2857d <= matchd2856d;
	-- d2858d
	sted2858d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2858d,
			Enable=>Enabled2858d,
			match=>matchd2858d,
			run=>run);

	Enabled2858d <= matchd2857d;
	-- d2859d
	sted2859d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2859d,
			Enable=>Enabled2859d,
			match=>matchd2859d,
			run=>run);

	Enabled2859d <= matchd2859d OR matchd2858d;
	-- d2860d
	sted2860d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2860d,
			Enable=>Enabled2860d,
			match=>matchd2860d,
			run=>run);

	Enabled2860d <= matchd2859d;
	-- d2861d
	sted2861d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2861d,
			Enable=>Enabled2861d,
			match=>matchd2861d,
			run=>run);

	Enabled2861d <= matchd2860d OR matchd2861d;
	-- d2862d
	sted2862d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2862d,
			Enable=>Enabled2862d,
			match=>matchd2862d,
			run=>run);

	Enabled2862d <= matchd2861d;
	-- d2863d
	sted2863d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2863d,
			Enable=>Enabled2863d,
			match=>matchd2863d,
			run=>run);

	Enabled2863d <= matchd2862d OR matchd2863d;
	-- d2864d
	sted2864d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2864d,
			Enable=>Enabled2864d,
			match=>matchd2864d,
			run=>run);

	Enabled2864d <= matchd2863d;
	-- d2865d
	sted2865d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2865d,
			Enable=>Enabled2865d,
			match=>matchd2865d,
			run=>run);

	Enabled2865d <= matchd2864d;
	-- d2866d
	sted2866d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2866d,
			Enable=>Enabled2866d,
			match=>matchd2866d,
			run=>run);

	Enabled2866d <= matchd2865d;
	-- d2867d
	sted2867d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2867d,
			Enable=>Enabled2867d,
			match=>matchd2867d,
			run=>run);

	Enabled2867d <= matchd2866d;
	-- d2868d
	sted2868d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2868d,
			Enable=>Enabled2868d,
			match=>matchd2868d,
			run=>run);

	Enabled2868d <= matchd2867d;
	-- d2870d
	sted2870d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2870d,
			Enable=>Enabled2870d,
			match=>matchd2870d,
			run=>run);

	-- d2871d
	sted2871d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2871d,
			Enable=>Enabled2871d,
			match=>matchd2871d,
			run=>run);

	Enabled2871d <= matchd2871d OR matchd2870d;
	-- d2872d
	sted2872d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2872d,
			Enable=>Enabled2872d,
			match=>matchd2872d,
			run=>run);

	Enabled2872d <= matchd2871d;
	-- d2873d
	sted2873d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2873d,
			Enable=>Enabled2873d,
			match=>matchd2873d,
			run=>run);

	Enabled2873d <= matchd2872d;
	-- d2874d
	sted2874d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2874d,
			Enable=>Enabled2874d,
			match=>matchd2874d,
			run=>run);

	Enabled2874d <= matchd2873d;
	-- d2875d
	sted2875d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2875d,
			Enable=>Enabled2875d,
			match=>matchd2875d,
			run=>run);

	Enabled2875d <= matchd2874d;
	-- d2876d
	sted2876d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2876d,
			Enable=>Enabled2876d,
			match=>matchd2876d,
			run=>run);

	Enabled2876d <= matchd2875d;
	-- d2877d
	sted2877d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2877d,
			Enable=>Enabled2877d,
			match=>matchd2877d,
			run=>run);

	Enabled2877d <= matchd2877d OR matchd2876d;
	-- d2878d
	sted2878d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2878d,
			Enable=>Enabled2878d,
			match=>matchd2878d,
			run=>run);

	Enabled2878d <= matchd2877d;
	-- d2879d
	sted2879d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2879d,
			Enable=>Enabled2879d,
			match=>matchd2879d,
			run=>run);

	Enabled2879d <= matchd2878d;
	-- d2880d
	sted2880d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2880d,
			Enable=>Enabled2880d,
			match=>matchd2880d,
			run=>run);

	Enabled2880d <= matchd2879d;
	-- d2881d
	sted2881d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2881d,
			Enable=>Enabled2881d,
			match=>matchd2881d,
			run=>run);

	Enabled2881d <= matchd2880d;
	-- d2882d
	sted2882d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2882d,
			Enable=>Enabled2882d,
			match=>matchd2882d,
			run=>run);

	reports(154) <= matchd2882d;
	Enabled2882d <= matchd2881d;
	-- d2883d
	sted2883d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2883d,
			Enable=>Enabled2883d,
			match=>matchd2883d,
			run=>run);

	-- d2884d
	sted2884d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2884d,
			Enable=>Enabled2884d,
			match=>matchd2884d,
			run=>run);

	Enabled2884d <= matchd2883d OR matchd2884d;
	-- d2885d
	sted2885d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2885d,
			Enable=>Enabled2885d,
			match=>matchd2885d,
			run=>run);

	Enabled2885d <= matchd2884d;
	-- d2886d
	sted2886d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2886d,
			Enable=>Enabled2886d,
			match=>matchd2886d,
			run=>run);

	Enabled2886d <= matchd2885d;
	-- d2887d
	sted2887d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2887d,
			Enable=>Enabled2887d,
			match=>matchd2887d,
			run=>run);

	Enabled2887d <= matchd2886d;
	-- d2888d
	sted2888d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2888d,
			Enable=>Enabled2888d,
			match=>matchd2888d,
			run=>run);

	Enabled2888d <= matchd2887d;
	-- d2889d
	sted2889d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2889d,
			Enable=>Enabled2889d,
			match=>matchd2889d,
			run=>run);

	Enabled2889d <= matchd2888d OR matchd2889d;
	-- d2890d
	sted2890d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2890d,
			Enable=>Enabled2890d,
			match=>matchd2890d,
			run=>run);

	Enabled2890d <= matchd2889d;
	-- d2891d
	sted2891d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2891d,
			Enable=>Enabled2891d,
			match=>matchd2891d,
			run=>run);

	Enabled2891d <= matchd2890d;
	-- d2892d
	sted2892d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2892d,
			Enable=>Enabled2892d,
			match=>matchd2892d,
			run=>run);

	Enabled2892d <= matchd2891d;
	-- d2893d
	sted2893d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2893d,
			Enable=>Enabled2893d,
			match=>matchd2893d,
			run=>run);

	Enabled2893d <= matchd2892d;
	-- d2894d
	sted2894d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2894d,
			Enable=>Enabled2894d,
			match=>matchd2894d,
			run=>run);

	Enabled2894d <= matchd2893d OR matchd2894d;
	-- d2895d
	sted2895d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2895d,
			Enable=>Enabled2895d,
			match=>matchd2895d,
			run=>run);

	Enabled2895d <= matchd2894d;
	-- d2896d
	sted2896d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2896d,
			Enable=>Enabled2896d,
			match=>matchd2896d,
			run=>run);

	Enabled2896d <= matchd2895d;
	-- d2897d
	sted2897d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2897d,
			Enable=>Enabled2897d,
			match=>matchd2897d,
			run=>run);

	Enabled2897d <= matchd2896d;
	-- d2898d
	sted2898d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2898d,
			Enable=>Enabled2898d,
			match=>matchd2898d,
			run=>run);

	Enabled2898d <= matchd2897d;
	-- d2899d
	sted2899d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2899d,
			Enable=>Enabled2899d,
			match=>matchd2899d,
			run=>run);

	reports(155) <= matchd2899d;
	Enabled2899d <= matchd2898d;
	-- d2900d
	sted2900d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2900d,
			Enable=>Enabled2900d,
			match=>matchd2900d,
			run=>run);

	-- d2901d
	sted2901d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2901d,
			Enable=>Enabled2901d,
			match=>matchd2901d,
			run=>run);

	Enabled2901d <= matchd2901d OR matchd2900d;
	-- d2902d
	sted2902d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2902d,
			Enable=>Enabled2902d,
			match=>matchd2902d,
			run=>run);

	Enabled2902d <= matchd2901d;
	-- d2903d
	sted2903d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2903d,
			Enable=>Enabled2903d,
			match=>matchd2903d,
			run=>run);

	Enabled2903d <= matchd2902d;
	-- d2904d
	sted2904d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2904d,
			Enable=>Enabled2904d,
			match=>matchd2904d,
			run=>run);

	Enabled2904d <= matchd2903d;
	-- d2905d
	sted2905d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2905d,
			Enable=>Enabled2905d,
			match=>matchd2905d,
			run=>run);

	Enabled2905d <= matchd2904d;
	-- d2906d
	sted2906d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2906d,
			Enable=>Enabled2906d,
			match=>matchd2906d,
			run=>run);

	Enabled2906d <= matchd2905d;
	-- d2907d
	sted2907d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2907d,
			Enable=>Enabled2907d,
			match=>matchd2907d,
			run=>run);

	Enabled2907d <= matchd2907d OR matchd2906d;
	-- d2908d
	sted2908d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2908d,
			Enable=>Enabled2908d,
			match=>matchd2908d,
			run=>run);

	Enabled2908d <= matchd2907d;
	-- d2909d
	sted2909d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2909d,
			Enable=>Enabled2909d,
			match=>matchd2909d,
			run=>run);

	Enabled2909d <= matchd2908d;
	-- d2910d
	sted2910d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2910d,
			Enable=>Enabled2910d,
			match=>matchd2910d,
			run=>run);

	Enabled2910d <= matchd2909d;
	-- d2911d
	sted2911d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2911d,
			Enable=>Enabled2911d,
			match=>matchd2911d,
			run=>run);

	Enabled2911d <= matchd2910d;
	-- d2912d
	sted2912d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2912d,
			Enable=>Enabled2912d,
			match=>matchd2912d,
			run=>run);

	reports(156) <= matchd2912d;
	Enabled2912d <= matchd2911d;
	-- d2913d
	sted2913d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2913d,
			Enable=>Enabled2913d,
			match=>matchd2913d,
			run=>run);

	-- d2914d
	sted2914d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2914d,
			Enable=>Enabled2914d,
			match=>matchd2914d,
			run=>run);

	Enabled2914d <= matchd2913d;
	-- d2915d
	sted2915d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2915d,
			Enable=>Enabled2915d,
			match=>matchd2915d,
			run=>run);

	Enabled2915d <= matchd2914d;
	-- d2916d
	sted2916d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2916d,
			Enable=>Enabled2916d,
			match=>matchd2916d,
			run=>run);

	Enabled2916d <= matchd2915d;
	-- d2917d
	sted2917d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2917d,
			Enable=>Enabled2917d,
			match=>matchd2917d,
			run=>run);

	Enabled2917d <= matchd2916d;
	-- d2918d
	sted2918d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2918d,
			Enable=>Enabled2918d,
			match=>matchd2918d,
			run=>run);

	Enabled2918d <= matchd2917d;
	-- d2919d
	sted2919d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2919d,
			Enable=>Enabled2919d,
			match=>matchd2919d,
			run=>run);

	Enabled2919d <= matchd2918d;
	-- d2920d
	sted2920d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2920d,
			Enable=>Enabled2920d,
			match=>matchd2920d,
			run=>run);

	Enabled2920d <= matchd2920d OR matchd2919d;
	-- d2921d
	sted2921d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2921d,
			Enable=>Enabled2921d,
			match=>matchd2921d,
			run=>run);

	Enabled2921d <= matchd2920d;
	-- d2922d
	sted2922d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2922d,
			Enable=>Enabled2922d,
			match=>matchd2922d,
			run=>run);

	Enabled2922d <= matchd2921d;
	-- d2923d
	sted2923d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2923d,
			Enable=>Enabled2923d,
			match=>matchd2923d,
			run=>run);

	Enabled2923d <= matchd2922d;
	-- d2924d
	sted2924d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2924d,
			Enable=>Enabled2924d,
			match=>matchd2924d,
			run=>run);

	reports(157) <= matchd2924d;
	Enabled2924d <= matchd2923d;
	-- d2925d
	sted2925d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2925d,
			Enable=>Enabled2925d,
			match=>matchd2925d,
			run=>run);

	-- d2926d
	sted2926d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2926d,
			Enable=>Enabled2926d,
			match=>matchd2926d,
			run=>run);

	Enabled2926d <= matchd2925d;
	-- d2927d
	sted2927d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2927d,
			Enable=>Enabled2927d,
			match=>matchd2927d,
			run=>run);

	Enabled2927d <= matchd2926d;
	-- d2928d
	sted2928d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2928d,
			Enable=>Enabled2928d,
			match=>matchd2928d,
			run=>run);

	Enabled2928d <= matchd2927d;
	-- d2929d
	sted2929d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2929d,
			Enable=>Enabled2929d,
			match=>matchd2929d,
			run=>run);

	Enabled2929d <= matchd2928d;
	-- d2930d
	sted2930d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2930d,
			Enable=>Enabled2930d,
			match=>matchd2930d,
			run=>run);

	Enabled2930d <= matchd2929d;
	-- d2931d
	sted2931d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2931d,
			Enable=>Enabled2931d,
			match=>matchd2931d,
			run=>run);

	Enabled2931d <= matchd2930d;
	-- d2932d
	sted2932d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2932d,
			Enable=>Enabled2932d,
			match=>matchd2932d,
			run=>run);

	Enabled2932d <= matchd2931d;
	-- d2933d
	sted2933d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2933d,
			Enable=>Enabled2933d,
			match=>matchd2933d,
			run=>run);

	Enabled2933d <= matchd2932d;
	-- d2934d
	sted2934d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2934d,
			Enable=>Enabled2934d,
			match=>matchd2934d,
			run=>run);

	Enabled2934d <= matchd2933d;
	-- d2935d
	sted2935d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2935d,
			Enable=>Enabled2935d,
			match=>matchd2935d,
			run=>run);

	Enabled2935d <= matchd2934d;
	-- d2936d
	sted2936d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2936d,
			Enable=>Enabled2936d,
			match=>matchd2936d,
			run=>run);

	Enabled2936d <= matchd2935d OR matchd2936d;
	-- d2937d
	sted2937d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2937d,
			Enable=>Enabled2937d,
			match=>matchd2937d,
			run=>run);

	Enabled2937d <= matchd2936d;
	-- d2938d
	sted2938d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2938d,
			Enable=>Enabled2938d,
			match=>matchd2938d,
			run=>run);

	Enabled2938d <= matchd2937d;
	-- d2939d
	sted2939d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2939d,
			Enable=>Enabled2939d,
			match=>matchd2939d,
			run=>run);

	Enabled2939d <= matchd2938d;
	-- d2940d
	sted2940d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2940d,
			Enable=>Enabled2940d,
			match=>matchd2940d,
			run=>run);

	Enabled2940d <= matchd2939d;
	-- d2941d
	sted2941d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2941d,
			Enable=>Enabled2941d,
			match=>matchd2941d,
			run=>run);

	reports(158) <= matchd2941d;
	Enabled2941d <= matchd2940d;
	-- d2942d
	sted2942d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2942d,
			Enable=>Enabled2942d,
			match=>matchd2942d,
			run=>run);

	-- d2943d
	sted2943d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2943d,
			Enable=>Enabled2943d,
			match=>matchd2943d,
			run=>run);

	Enabled2943d <= matchd2942d;
	-- d2944d
	sted2944d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2944d,
			Enable=>Enabled2944d,
			match=>matchd2944d,
			run=>run);

	Enabled2944d <= matchd2943d;
	-- d2945d
	sted2945d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2945d,
			Enable=>Enabled2945d,
			match=>matchd2945d,
			run=>run);

	Enabled2945d <= matchd2944d;
	-- d2946d
	sted2946d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2946d,
			Enable=>Enabled2946d,
			match=>matchd2946d,
			run=>run);

	Enabled2946d <= matchd2945d;
	-- d2947d
	sted2947d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2947d,
			Enable=>Enabled2947d,
			match=>matchd2947d,
			run=>run);

	Enabled2947d <= matchd2946d;
	-- d2948d
	sted2948d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2948d,
			Enable=>Enabled2948d,
			match=>matchd2948d,
			run=>run);

	Enabled2948d <= matchd2947d;
	-- d2949d
	sted2949d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2949d,
			Enable=>Enabled2949d,
			match=>matchd2949d,
			run=>run);

	Enabled2949d <= matchd2948d;
	-- d2950d
	sted2950d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2950d,
			Enable=>Enabled2950d,
			match=>matchd2950d,
			run=>run);

	Enabled2950d <= matchd2949d;
	-- d2951d
	sted2951d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2951d,
			Enable=>Enabled2951d,
			match=>matchd2951d,
			run=>run);

	Enabled2951d <= matchd2950d;
	-- d2952d
	sted2952d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2952d,
			Enable=>Enabled2952d,
			match=>matchd2952d,
			run=>run);

	Enabled2952d <= matchd2952d OR matchd2951d;
	-- d2953d
	sted2953d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2953d,
			Enable=>Enabled2953d,
			match=>matchd2953d,
			run=>run);

	Enabled2953d <= matchd2952d;
	-- d2954d
	sted2954d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2954d,
			Enable=>Enabled2954d,
			match=>matchd2954d,
			run=>run);

	Enabled2954d <= matchd2953d;
	-- d2955d
	sted2955d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2955d,
			Enable=>Enabled2955d,
			match=>matchd2955d,
			run=>run);

	Enabled2955d <= matchd2954d;
	-- d2956d
	sted2956d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2956d,
			Enable=>Enabled2956d,
			match=>matchd2956d,
			run=>run);

	reports(159) <= matchd2956d;
	Enabled2956d <= matchd2955d;
	-- d2957d
	sted2957d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2957d,
			Enable=>Enabled2957d,
			match=>matchd2957d,
			run=>run);

	-- d2958d
	sted2958d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2958d,
			Enable=>Enabled2958d,
			match=>matchd2958d,
			run=>run);

	Enabled2958d <= matchd2958d OR matchd2957d;
	-- d2959d
	sted2959d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2959d,
			Enable=>Enabled2959d,
			match=>matchd2959d,
			run=>run);

	Enabled2959d <= matchd2958d;
	-- d2960d
	sted2960d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2960d,
			Enable=>Enabled2960d,
			match=>matchd2960d,
			run=>run);

	Enabled2960d <= matchd2959d;
	-- d2961d
	sted2961d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2961d,
			Enable=>Enabled2961d,
			match=>matchd2961d,
			run=>run);

	Enabled2961d <= matchd2960d;
	-- d2962d
	sted2962d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2962d,
			Enable=>Enabled2962d,
			match=>matchd2962d,
			run=>run);

	Enabled2962d <= matchd2961d;
	-- d2963d
	sted2963d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2963d,
			Enable=>Enabled2963d,
			match=>matchd2963d,
			run=>run);

	Enabled2963d <= matchd2962d OR matchd2963d;
	-- d2964d
	sted2964d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2964d,
			Enable=>Enabled2964d,
			match=>matchd2964d,
			run=>run);

	Enabled2964d <= matchd2963d;
	-- d2965d
	sted2965d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2965d,
			Enable=>Enabled2965d,
			match=>matchd2965d,
			run=>run);

	Enabled2965d <= matchd2964d;
	-- d2966d
	sted2966d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2966d,
			Enable=>Enabled2966d,
			match=>matchd2966d,
			run=>run);

	Enabled2966d <= matchd2965d;
	-- d2967d
	sted2967d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2967d,
			Enable=>Enabled2967d,
			match=>matchd2967d,
			run=>run);

	reports(160) <= matchd2967d;
	Enabled2967d <= matchd2966d;
	-- d2968d
	sted2968d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2968d,
			Enable=>Enabled2968d,
			match=>matchd2968d,
			run=>run);

	-- d2969d
	sted2969d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2969d,
			Enable=>Enabled2969d,
			match=>matchd2969d,
			run=>run);

	Enabled2969d <= matchd2968d OR matchd2969d;
	-- d2970d
	sted2970d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2970d,
			Enable=>Enabled2970d,
			match=>matchd2970d,
			run=>run);

	Enabled2970d <= matchd2969d;
	-- d2971d
	sted2971d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2971d,
			Enable=>Enabled2971d,
			match=>matchd2971d,
			run=>run);

	Enabled2971d <= matchd2970d;
	-- d2972d
	sted2972d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2972d,
			Enable=>Enabled2972d,
			match=>matchd2972d,
			run=>run);

	Enabled2972d <= matchd2971d;
	-- d2973d
	sted2973d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2973d,
			Enable=>Enabled2973d,
			match=>matchd2973d,
			run=>run);

	Enabled2973d <= matchd2972d;
	-- d2974d
	sted2974d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2974d,
			Enable=>Enabled2974d,
			match=>matchd2974d,
			run=>run);

	Enabled2974d <= matchd2973d OR matchd2974d;
	-- d2975d
	sted2975d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2975d,
			Enable=>Enabled2975d,
			match=>matchd2975d,
			run=>run);

	Enabled2975d <= matchd2974d;
	-- d2976d
	sted2976d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2976d,
			Enable=>Enabled2976d,
			match=>matchd2976d,
			run=>run);

	Enabled2976d <= matchd2975d;
	-- d2977d
	sted2977d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2977d,
			Enable=>Enabled2977d,
			match=>matchd2977d,
			run=>run);

	Enabled2977d <= matchd2976d;
	-- d2978d
	sted2978d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2978d,
			Enable=>Enabled2978d,
			match=>matchd2978d,
			run=>run);

	Enabled2978d <= matchd2977d;
	-- d2979d
	sted2979d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2979d,
			Enable=>Enabled2979d,
			match=>matchd2979d,
			run=>run);

	reports(161) <= matchd2979d;
	Enabled2979d <= matchd2978d;
	-- d2980d
	sted2980d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2980d,
			Enable=>Enabled2980d,
			match=>matchd2980d,
			run=>run);

	-- d2981d
	sted2981d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2981d,
			Enable=>Enabled2981d,
			match=>matchd2981d,
			run=>run);

	Enabled2981d <= matchd2981d OR matchd2980d;
	-- d2982d
	sted2982d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2982d,
			Enable=>Enabled2982d,
			match=>matchd2982d,
			run=>run);

	Enabled2982d <= matchd2981d;
	-- d2983d
	sted2983d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2983d,
			Enable=>Enabled2983d,
			match=>matchd2983d,
			run=>run);

	Enabled2983d <= matchd2982d;
	-- d2984d
	sted2984d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2984d,
			Enable=>Enabled2984d,
			match=>matchd2984d,
			run=>run);

	Enabled2984d <= matchd2983d;
	-- d2985d
	sted2985d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2985d,
			Enable=>Enabled2985d,
			match=>matchd2985d,
			run=>run);

	Enabled2985d <= matchd2984d;
	-- d2986d
	sted2986d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2986d,
			Enable=>Enabled2986d,
			match=>matchd2986d,
			run=>run);

	Enabled2986d <= matchd2985d;
	-- d2987d
	sted2987d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2987d,
			Enable=>Enabled2987d,
			match=>matchd2987d,
			run=>run);

	Enabled2987d <= matchd2986d;
	-- d2988d
	sted2988d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2988d,
			Enable=>Enabled2988d,
			match=>matchd2988d,
			run=>run);

	Enabled2988d <= matchd2988d OR matchd2987d;
	-- d2989d
	sted2989d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2989d,
			Enable=>Enabled2989d,
			match=>matchd2989d,
			run=>run);

	Enabled2989d <= matchd2988d;
	-- d2990d
	sted2990d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2990d,
			Enable=>Enabled2990d,
			match=>matchd2990d,
			run=>run);

	Enabled2990d <= matchd2989d;
	-- d2991d
	sted2991d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2991d,
			Enable=>Enabled2991d,
			match=>matchd2991d,
			run=>run);

	Enabled2991d <= matchd2990d;
	-- d2992d
	sted2992d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2992d,
			Enable=>Enabled2992d,
			match=>matchd2992d,
			run=>run);

	Enabled2992d <= matchd2991d;
	-- d2993d
	sted2993d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2993d,
			Enable=>Enabled2993d,
			match=>matchd2993d,
			run=>run);

	reports(162) <= matchd2993d;
	Enabled2993d <= matchd2992d;
	-- d2994d
	sted2994d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2994d,
			Enable=>Enabled2994d,
			match=>matchd2994d,
			run=>run);

	-- d2995d
	sted2995d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2995d,
			Enable=>Enabled2995d,
			match=>matchd2995d,
			run=>run);

	Enabled2995d <= matchd2994d;
	-- d2996d
	sted2996d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2996d,
			Enable=>Enabled2996d,
			match=>matchd2996d,
			run=>run);

	Enabled2996d <= matchd2995d;
	-- d2997d
	sted2997d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2997d,
			Enable=>Enabled2997d,
			match=>matchd2997d,
			run=>run);

	Enabled2997d <= matchd2996d;
	-- d2998d
	sted2998d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2998d,
			Enable=>Enabled2998d,
			match=>matchd2998d,
			run=>run);

	Enabled2998d <= matchd2997d;
	-- d2999d
	sted2999d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord2999d,
			Enable=>Enabled2999d,
			match=>matchd2999d,
			run=>run);

	Enabled2999d <= matchd2998d;
	-- d3000d
	sted3000d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3000d,
			Enable=>Enabled3000d,
			match=>matchd3000d,
			run=>run);

	Enabled3000d <= matchd2999d;
	-- d3001d
	sted3001d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3001d,
			Enable=>Enabled3001d,
			match=>matchd3001d,
			run=>run);

	Enabled3001d <= matchd3000d;
	-- d3002d
	sted3002d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3002d,
			Enable=>Enabled3002d,
			match=>matchd3002d,
			run=>run);

	Enabled3002d <= matchd3001d OR matchd3002d;
	-- d3003d
	sted3003d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3003d,
			Enable=>Enabled3003d,
			match=>matchd3003d,
			run=>run);

	Enabled3003d <= matchd3002d;
	-- d3004d
	sted3004d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3004d,
			Enable=>Enabled3004d,
			match=>matchd3004d,
			run=>run);

	Enabled3004d <= matchd3003d;
	-- d3005d
	sted3005d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3005d,
			Enable=>Enabled3005d,
			match=>matchd3005d,
			run=>run);

	Enabled3005d <= matchd3004d;
	-- d3006d
	sted3006d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3006d,
			Enable=>Enabled3006d,
			match=>matchd3006d,
			run=>run);

	Enabled3006d <= matchd3005d;
	-- d3007d
	sted3007d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3007d,
			Enable=>Enabled3007d,
			match=>matchd3007d,
			run=>run);

	reports(163) <= matchd3007d;
	Enabled3007d <= matchd3006d;
	-- d3008d
	sted3008d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3008d,
			Enable=>Enabled3008d,
			match=>matchd3008d,
			run=>run);

	-- d3009d
	sted3009d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3009d,
			Enable=>Enabled3009d,
			match=>matchd3009d,
			run=>run);

	Enabled3009d <= matchd3008d OR matchd3009d;
	-- d3010d
	sted3010d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3010d,
			Enable=>Enabled3010d,
			match=>matchd3010d,
			run=>run);

	Enabled3010d <= matchd3009d;
	-- d3011d
	sted3011d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3011d,
			Enable=>Enabled3011d,
			match=>matchd3011d,
			run=>run);

	Enabled3011d <= matchd3010d;
	-- d3012d
	sted3012d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3012d,
			Enable=>Enabled3012d,
			match=>matchd3012d,
			run=>run);

	Enabled3012d <= matchd3011d;
	-- d3013d
	sted3013d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3013d,
			Enable=>Enabled3013d,
			match=>matchd3013d,
			run=>run);

	Enabled3013d <= matchd3012d;
	-- d3014d
	sted3014d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3014d,
			Enable=>Enabled3014d,
			match=>matchd3014d,
			run=>run);

	Enabled3014d <= matchd3013d;
	-- d3015d
	sted3015d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3015d,
			Enable=>Enabled3015d,
			match=>matchd3015d,
			run=>run);

	Enabled3015d <= matchd3014d;
	-- d3016d
	sted3016d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3016d,
			Enable=>Enabled3016d,
			match=>matchd3016d,
			run=>run);

	Enabled3016d <= matchd3015d;
	-- d3017d
	sted3017d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3017d,
			Enable=>Enabled3017d,
			match=>matchd3017d,
			run=>run);

	Enabled3017d <= matchd3016d;
	-- d3018d
	sted3018d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3018d,
			Enable=>Enabled3018d,
			match=>matchd3018d,
			run=>run);

	Enabled3018d <= matchd3017d;
	-- d3019d
	sted3019d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3019d,
			Enable=>Enabled3019d,
			match=>matchd3019d,
			run=>run);

	Enabled3019d <= matchd3018d;
	-- d3020d
	sted3020d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3020d,
			Enable=>Enabled3020d,
			match=>matchd3020d,
			run=>run);

	Enabled3020d <= matchd3019d;
	-- d3021d
	sted3021d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3021d,
			Enable=>Enabled3021d,
			match=>matchd3021d,
			run=>run);

	Enabled3021d <= matchd3020d;
	-- d3022d
	sted3022d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3022d,
			Enable=>Enabled3022d,
			match=>matchd3022d,
			run=>run);

	Enabled3022d <= matchd3021d;
	-- d3023d
	sted3023d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3023d,
			Enable=>Enabled3023d,
			match=>matchd3023d,
			run=>run);

	reports(164) <= matchd3023d;
	Enabled3023d <= matchd3022d;
	-- d3024d
	sted3024d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3024d,
			Enable=>Enabled3024d,
			match=>matchd3024d,
			run=>run);

	-- d3025d
	sted3025d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3025d,
			Enable=>Enabled3025d,
			match=>matchd3025d,
			run=>run);

	Enabled3025d <= matchd3024d OR matchd3025d;
	-- d3026d
	sted3026d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3026d,
			Enable=>Enabled3026d,
			match=>matchd3026d,
			run=>run);

	Enabled3026d <= matchd3025d;
	-- d3027d
	sted3027d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3027d,
			Enable=>Enabled3027d,
			match=>matchd3027d,
			run=>run);

	Enabled3027d <= matchd3026d;
	-- d3028d
	sted3028d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3028d,
			Enable=>Enabled3028d,
			match=>matchd3028d,
			run=>run);

	Enabled3028d <= matchd3027d;
	-- d3029d
	sted3029d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3029d,
			Enable=>Enabled3029d,
			match=>matchd3029d,
			run=>run);

	Enabled3029d <= matchd3028d;
	-- d3030d
	sted3030d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3030d,
			Enable=>Enabled3030d,
			match=>matchd3030d,
			run=>run);

	Enabled3030d <= matchd3029d;
	-- d3031d
	sted3031d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3031d,
			Enable=>Enabled3031d,
			match=>matchd3031d,
			run=>run);

	Enabled3031d <= matchd3030d;
	-- d3032d
	sted3032d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3032d,
			Enable=>Enabled3032d,
			match=>matchd3032d,
			run=>run);

	Enabled3032d <= matchd3031d;
	-- d3033d
	sted3033d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3033d,
			Enable=>Enabled3033d,
			match=>matchd3033d,
			run=>run);

	Enabled3033d <= matchd3032d;
	-- d3034d
	sted3034d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3034d,
			Enable=>Enabled3034d,
			match=>matchd3034d,
			run=>run);

	Enabled3034d <= matchd3033d;
	-- d3035d
	sted3035d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3035d,
			Enable=>Enabled3035d,
			match=>matchd3035d,
			run=>run);

	Enabled3035d <= matchd3034d OR matchd3035d;
	-- d3036d
	sted3036d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3036d,
			Enable=>Enabled3036d,
			match=>matchd3036d,
			run=>run);

	Enabled3036d <= matchd3035d;
	-- d3037d
	sted3037d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3037d,
			Enable=>Enabled3037d,
			match=>matchd3037d,
			run=>run);

	Enabled3037d <= matchd3037d OR matchd3036d;
	-- d3038d
	sted3038d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3038d,
			Enable=>Enabled3038d,
			match=>matchd3038d,
			run=>run);

	Enabled3038d <= matchd3037d;
	-- d3039d
	sted3039d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3039d,
			Enable=>Enabled3039d,
			match=>matchd3039d,
			run=>run);

	Enabled3039d <= matchd3038d OR matchd3039d;
	-- d3040d
	sted3040d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3040d,
			Enable=>Enabled3040d,
			match=>matchd3040d,
			run=>run);

	Enabled3040d <= matchd3039d;
	-- d3041d
	sted3041d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3041d,
			Enable=>Enabled3041d,
			match=>matchd3041d,
			run=>run);

	-- d3042d
	sted3042d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3042d,
			Enable=>Enabled3042d,
			match=>matchd3042d,
			run=>run);

	Enabled3042d <= matchd3042d OR matchd3041d;
	-- d3043d
	sted3043d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3043d,
			Enable=>Enabled3043d,
			match=>matchd3043d,
			run=>run);

	Enabled3043d <= matchd3042d;
	-- d3044d
	sted3044d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3044d,
			Enable=>Enabled3044d,
			match=>matchd3044d,
			run=>run);

	Enabled3044d <= matchd3043d;
	-- d3045d
	sted3045d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3045d,
			Enable=>Enabled3045d,
			match=>matchd3045d,
			run=>run);

	Enabled3045d <= matchd3044d;
	-- d3046d
	sted3046d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3046d,
			Enable=>Enabled3046d,
			match=>matchd3046d,
			run=>run);

	Enabled3046d <= matchd3045d;
	-- d3047d
	sted3047d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3047d,
			Enable=>Enabled3047d,
			match=>matchd3047d,
			run=>run);

	Enabled3047d <= matchd3047d OR matchd3046d;
	-- d3048d
	sted3048d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3048d,
			Enable=>Enabled3048d,
			match=>matchd3048d,
			run=>run);

	Enabled3048d <= matchd3047d;
	-- d3049d
	sted3049d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3049d,
			Enable=>Enabled3049d,
			match=>matchd3049d,
			run=>run);

	Enabled3049d <= matchd3049d OR matchd3048d;
	-- d3050d
	sted3050d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3050d,
			Enable=>Enabled3050d,
			match=>matchd3050d,
			run=>run);

	Enabled3050d <= matchd3049d;
	-- d3051d
	sted3051d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3051d,
			Enable=>Enabled3051d,
			match=>matchd3051d,
			run=>run);

	Enabled3051d <= matchd3050d;
	-- d3052d
	sted3052d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3052d,
			Enable=>Enabled3052d,
			match=>matchd3052d,
			run=>run);

	Enabled3052d <= matchd3051d;
	-- d3053d
	sted3053d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3053d,
			Enable=>Enabled3053d,
			match=>matchd3053d,
			run=>run);

	Enabled3053d <= matchd3052d;
	-- d3054d
	sted3054d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3054d,
			Enable=>Enabled3054d,
			match=>matchd3054d,
			run=>run);

	Enabled3054d <= matchd3053d;
	-- d3055d
	sted3055d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3055d,
			Enable=>Enabled3055d,
			match=>matchd3055d,
			run=>run);

	Enabled3055d <= matchd3054d;
	-- d3056d
	sted3056d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3056d,
			Enable=>Enabled3056d,
			match=>matchd3056d,
			run=>run);

	Enabled3056d <= matchd3055d OR matchd3056d;
	-- d3057d
	sted3057d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3057d,
			Enable=>Enabled3057d,
			match=>matchd3057d,
			run=>run);

	Enabled3057d <= matchd3056d;
	-- d3059d
	sted3059d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3059d,
			Enable=>Enabled3059d,
			match=>matchd3059d,
			run=>run);

	-- d3060d
	sted3060d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3060d,
			Enable=>Enabled3060d,
			match=>matchd3060d,
			run=>run);

	Enabled3060d <= matchd3059d OR matchd3060d;
	-- d3061d
	sted3061d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3061d,
			Enable=>Enabled3061d,
			match=>matchd3061d,
			run=>run);

	Enabled3061d <= matchd3060d;
	-- d3062d
	sted3062d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3062d,
			Enable=>Enabled3062d,
			match=>matchd3062d,
			run=>run);

	Enabled3062d <= matchd3061d;
	-- d3063d
	sted3063d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3063d,
			Enable=>Enabled3063d,
			match=>matchd3063d,
			run=>run);

	Enabled3063d <= matchd3062d;
	-- d3064d
	sted3064d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3064d,
			Enable=>Enabled3064d,
			match=>matchd3064d,
			run=>run);

	Enabled3064d <= matchd3063d;
	-- d3065d
	sted3065d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3065d,
			Enable=>Enabled3065d,
			match=>matchd3065d,
			run=>run);

	Enabled3065d <= matchd3064d OR matchd3065d;
	-- d3066d
	sted3066d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3066d,
			Enable=>Enabled3066d,
			match=>matchd3066d,
			run=>run);

	Enabled3066d <= matchd3065d;
	-- d3067d
	sted3067d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3067d,
			Enable=>Enabled3067d,
			match=>matchd3067d,
			run=>run);

	Enabled3067d <= matchd3066d OR matchd3067d;
	-- d3068d
	sted3068d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3068d,
			Enable=>Enabled3068d,
			match=>matchd3068d,
			run=>run);

	Enabled3068d <= matchd3067d;
	-- d3069d
	sted3069d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3069d,
			Enable=>Enabled3069d,
			match=>matchd3069d,
			run=>run);

	Enabled3069d <= matchd3068d OR matchd3069d;
	-- d3070d
	sted3070d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3070d,
			Enable=>Enabled3070d,
			match=>matchd3070d,
			run=>run);

	Enabled3070d <= matchd3069d;
	-- d3071d
	sted3071d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3071d,
			Enable=>Enabled3071d,
			match=>matchd3071d,
			run=>run);

	Enabled3071d <= matchd3070d OR matchd3071d;
	-- d3072d
	sted3072d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3072d,
			Enable=>Enabled3072d,
			match=>matchd3072d,
			run=>run);

	Enabled3072d <= matchd3071d;
	-- d3073d
	sted3073d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3073d,
			Enable=>Enabled3073d,
			match=>matchd3073d,
			run=>run);

	Enabled3073d <= matchd3072d OR matchd3073d;
	-- d3074d
	sted3074d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3074d,
			Enable=>Enabled3074d,
			match=>matchd3074d,
			run=>run);

	Enabled3074d <= matchd3073d;
	-- d3075d
	sted3075d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3075d,
			Enable=>Enabled3075d,
			match=>matchd3075d,
			run=>run);

	Enabled3075d <= matchd3074d;
	-- d3076d
	sted3076d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3076d,
			Enable=>Enabled3076d,
			match=>matchd3076d,
			run=>run);

	Enabled3076d <= matchd3075d;
	-- d3077d
	sted3077d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3077d,
			Enable=>Enabled3077d,
			match=>matchd3077d,
			run=>run);

	Enabled3077d <= matchd3076d;
	-- d3078d
	sted3078d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3078d,
			Enable=>Enabled3078d,
			match=>matchd3078d,
			run=>run);

	-- d3079d
	sted3079d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3079d,
			Enable=>Enabled3079d,
			match=>matchd3079d,
			run=>run);

	Enabled3079d <= matchd3078d OR matchd3079d;
	-- d3080d
	sted3080d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3080d,
			Enable=>Enabled3080d,
			match=>matchd3080d,
			run=>run);

	Enabled3080d <= matchd3079d;
	-- d3081d
	sted3081d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3081d,
			Enable=>Enabled3081d,
			match=>matchd3081d,
			run=>run);

	Enabled3081d <= matchd3080d OR matchd3081d;
	-- d3082d
	sted3082d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3082d,
			Enable=>Enabled3082d,
			match=>matchd3082d,
			run=>run);

	Enabled3082d <= matchd3081d;
	-- d3083d
	sted3083d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3083d,
			Enable=>Enabled3083d,
			match=>matchd3083d,
			run=>run);

	Enabled3083d <= matchd3082d OR matchd3083d;
	-- d3084d
	sted3084d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3084d,
			Enable=>Enabled3084d,
			match=>matchd3084d,
			run=>run);

	Enabled3084d <= matchd3083d;
	-- d3085d
	sted3085d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3085d,
			Enable=>Enabled3085d,
			match=>matchd3085d,
			run=>run);

	Enabled3085d <= matchd3084d;
	-- d3086d
	sted3086d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3086d,
			Enable=>Enabled3086d,
			match=>matchd3086d,
			run=>run);

	Enabled3086d <= matchd3085d;
	-- d3087d
	sted3087d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3087d,
			Enable=>Enabled3087d,
			match=>matchd3087d,
			run=>run);

	Enabled3087d <= matchd3086d;
	-- d3088d
	sted3088d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3088d,
			Enable=>Enabled3088d,
			match=>matchd3088d,
			run=>run);

	Enabled3088d <= matchd3087d OR matchd3088d;
	-- d3089d
	sted3089d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3089d,
			Enable=>Enabled3089d,
			match=>matchd3089d,
			run=>run);

	Enabled3089d <= matchd3088d;
	-- d3090d
	sted3090d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3090d,
			Enable=>Enabled3090d,
			match=>matchd3090d,
			run=>run);

	Enabled3090d <= matchd3090d OR matchd3089d;
	-- d3091d
	sted3091d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3091d,
			Enable=>Enabled3091d,
			match=>matchd3091d,
			run=>run);

	Enabled3091d <= matchd3090d;
	-- d3092d
	sted3092d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3092d,
			Enable=>Enabled3092d,
			match=>matchd3092d,
			run=>run);

	Enabled3092d <= matchd3091d OR matchd3092d;
	-- d3093d
	sted3093d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3093d,
			Enable=>Enabled3093d,
			match=>matchd3093d,
			run=>run);

	Enabled3093d <= matchd3092d;
	-- d3094d
	sted3094d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3094d,
			Enable=>Enabled3094d,
			match=>matchd3094d,
			run=>run);

	Enabled3094d <= matchd3093d;
	-- d3095d
	sted3095d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3095d,
			Enable=>Enabled3095d,
			match=>matchd3095d,
			run=>run);

	Enabled3095d <= matchd3094d;
	-- d3096d
	sted3096d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3096d,
			Enable=>Enabled3096d,
			match=>matchd3096d,
			run=>run);

	Enabled3096d <= matchd3095d;
	-- d3097d
	sted3097d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3097d,
			Enable=>Enabled3097d,
			match=>matchd3097d,
			run=>run);

	-- d3098d
	sted3098d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3098d,
			Enable=>Enabled3098d,
			match=>matchd3098d,
			run=>run);

	Enabled3098d <= matchd3098d OR matchd3097d;
	-- d3099d
	sted3099d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3099d,
			Enable=>Enabled3099d,
			match=>matchd3099d,
			run=>run);

	Enabled3099d <= matchd3098d;
	-- d3100d
	sted3100d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3100d,
			Enable=>Enabled3100d,
			match=>matchd3100d,
			run=>run);

	Enabled3100d <= matchd3099d OR matchd3100d;
	-- d3101d
	sted3101d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3101d,
			Enable=>Enabled3101d,
			match=>matchd3101d,
			run=>run);

	Enabled3101d <= matchd3100d;
	-- d3102d
	sted3102d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3102d,
			Enable=>Enabled3102d,
			match=>matchd3102d,
			run=>run);

	Enabled3102d <= matchd3101d OR matchd3102d;
	-- d3103d
	sted3103d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3103d,
			Enable=>Enabled3103d,
			match=>matchd3103d,
			run=>run);

	Enabled3103d <= matchd3102d;
	-- d3104d
	sted3104d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3104d,
			Enable=>Enabled3104d,
			match=>matchd3104d,
			run=>run);

	Enabled3104d <= matchd3104d OR matchd3103d;
	-- d3105d
	sted3105d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3105d,
			Enable=>Enabled3105d,
			match=>matchd3105d,
			run=>run);

	Enabled3105d <= matchd3104d;
	-- d3106d
	sted3106d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3106d,
			Enable=>Enabled3106d,
			match=>matchd3106d,
			run=>run);

	Enabled3106d <= matchd3105d OR matchd3106d;
	-- d3107d
	sted3107d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3107d,
			Enable=>Enabled3107d,
			match=>matchd3107d,
			run=>run);

	Enabled3107d <= matchd3106d;
	-- d3108d
	sted3108d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3108d,
			Enable=>Enabled3108d,
			match=>matchd3108d,
			run=>run);

	Enabled3108d <= matchd3107d;
	-- d3109d
	sted3109d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3109d,
			Enable=>Enabled3109d,
			match=>matchd3109d,
			run=>run);

	Enabled3109d <= matchd3108d;
	-- d3110d
	sted3110d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3110d,
			Enable=>Enabled3110d,
			match=>matchd3110d,
			run=>run);

	Enabled3110d <= matchd3109d;
	-- d3111d
	sted3111d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3111d,
			Enable=>Enabled3111d,
			match=>matchd3111d,
			run=>run);

	Enabled3111d <= matchd3111d OR matchd3110d;
	-- d3112d
	sted3112d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3112d,
			Enable=>Enabled3112d,
			match=>matchd3112d,
			run=>run);

	Enabled3112d <= matchd3111d;
	-- d3113d
	sted3113d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3113d,
			Enable=>Enabled3113d,
			match=>matchd3113d,
			run=>run);

	Enabled3113d <= matchd3112d;
	-- d3114d
	sted3114d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3114d,
			Enable=>Enabled3114d,
			match=>matchd3114d,
			run=>run);

	Enabled3114d <= matchd3113d;
	-- d3115d
	sted3115d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3115d,
			Enable=>Enabled3115d,
			match=>matchd3115d,
			run=>run);

	Enabled3115d <= matchd3114d;
	-- d3117d
	sted3117d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3117d,
			Enable=>Enabled3117d,
			match=>matchd3117d,
			run=>run);

	-- d3118d
	sted3118d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3118d,
			Enable=>Enabled3118d,
			match=>matchd3118d,
			run=>run);

	Enabled3118d <= matchd3118d OR matchd3117d;
	-- d3119d
	sted3119d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3119d,
			Enable=>Enabled3119d,
			match=>matchd3119d,
			run=>run);

	Enabled3119d <= matchd3118d;
	-- d3120d
	sted3120d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3120d,
			Enable=>Enabled3120d,
			match=>matchd3120d,
			run=>run);

	Enabled3120d <= matchd3119d;
	-- d3121d
	sted3121d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3121d,
			Enable=>Enabled3121d,
			match=>matchd3121d,
			run=>run);

	Enabled3121d <= matchd3120d;
	-- d3122d
	sted3122d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3122d,
			Enable=>Enabled3122d,
			match=>matchd3122d,
			run=>run);

	Enabled3122d <= matchd3121d;
	-- d3123d
	sted3123d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3123d,
			Enable=>Enabled3123d,
			match=>matchd3123d,
			run=>run);

	Enabled3123d <= matchd3122d;
	-- d3124d
	sted3124d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3124d,
			Enable=>Enabled3124d,
			match=>matchd3124d,
			run=>run);

	Enabled3124d <= matchd3123d;
	-- d3125d
	sted3125d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3125d,
			Enable=>Enabled3125d,
			match=>matchd3125d,
			run=>run);

	Enabled3125d <= matchd3124d OR matchd3125d;
	-- d3126d
	sted3126d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3126d,
			Enable=>Enabled3126d,
			match=>matchd3126d,
			run=>run);

	Enabled3126d <= matchd3125d;
	-- d3127d
	sted3127d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3127d,
			Enable=>Enabled3127d,
			match=>matchd3127d,
			run=>run);

	Enabled3127d <= matchd3126d;
	-- d3128d
	sted3128d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3128d,
			Enable=>Enabled3128d,
			match=>matchd3128d,
			run=>run);

	Enabled3128d <= matchd3127d;
	-- d3129d
	sted3129d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3129d,
			Enable=>Enabled3129d,
			match=>matchd3129d,
			run=>run);

	Enabled3129d <= matchd3128d;
	-- d3130d
	sted3130d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3130d,
			Enable=>Enabled3130d,
			match=>matchd3130d,
			run=>run);

	reports(165) <= matchd3130d;
	Enabled3130d <= matchd3129d;
	-- d3131d
	sted3131d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3131d,
			Enable=>Enabled3131d,
			match=>matchd3131d,
			run=>run);

	-- d3132d
	sted3132d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3132d,
			Enable=>Enabled3132d,
			match=>matchd3132d,
			run=>run);

	Enabled3132d <= matchd3131d OR matchd3132d;
	-- d3133d
	sted3133d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3133d,
			Enable=>Enabled3133d,
			match=>matchd3133d,
			run=>run);

	Enabled3133d <= matchd3132d;
	-- d3134d
	sted3134d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3134d,
			Enable=>Enabled3134d,
			match=>matchd3134d,
			run=>run);

	Enabled3134d <= matchd3133d;
	-- d3135d
	sted3135d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3135d,
			Enable=>Enabled3135d,
			match=>matchd3135d,
			run=>run);

	Enabled3135d <= matchd3134d;
	-- d3136d
	sted3136d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3136d,
			Enable=>Enabled3136d,
			match=>matchd3136d,
			run=>run);

	Enabled3136d <= matchd3135d;
	-- d3137d
	sted3137d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3137d,
			Enable=>Enabled3137d,
			match=>matchd3137d,
			run=>run);

	Enabled3137d <= matchd3136d;
	-- d3138d
	sted3138d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3138d,
			Enable=>Enabled3138d,
			match=>matchd3138d,
			run=>run);

	Enabled3138d <= matchd3137d OR matchd3138d;
	-- d3139d
	sted3139d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3139d,
			Enable=>Enabled3139d,
			match=>matchd3139d,
			run=>run);

	Enabled3139d <= matchd3138d;
	-- d3140d
	sted3140d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3140d,
			Enable=>Enabled3140d,
			match=>matchd3140d,
			run=>run);

	Enabled3140d <= matchd3139d;
	-- d3141d
	sted3141d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3141d,
			Enable=>Enabled3141d,
			match=>matchd3141d,
			run=>run);

	Enabled3141d <= matchd3140d;
	-- d3142d
	sted3142d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3142d,
			Enable=>Enabled3142d,
			match=>matchd3142d,
			run=>run);

	Enabled3142d <= matchd3141d;
	-- d3143d
	sted3143d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3143d,
			Enable=>Enabled3143d,
			match=>matchd3143d,
			run=>run);

	Enabled3143d <= matchd3142d;
	-- d3144d
	sted3144d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3144d,
			Enable=>Enabled3144d,
			match=>matchd3144d,
			run=>run);

	Enabled3144d <= matchd3143d OR matchd3144d;
	-- d3145d
	sted3145d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3145d,
			Enable=>Enabled3145d,
			match=>matchd3145d,
			run=>run);

	Enabled3145d <= matchd3144d;
	-- d3146d
	sted3146d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3146d,
			Enable=>Enabled3146d,
			match=>matchd3146d,
			run=>run);

	Enabled3146d <= matchd3145d;
	-- d3147d
	sted3147d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3147d,
			Enable=>Enabled3147d,
			match=>matchd3147d,
			run=>run);

	Enabled3147d <= matchd3146d;
	-- d3148d
	sted3148d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3148d,
			Enable=>Enabled3148d,
			match=>matchd3148d,
			run=>run);

	Enabled3148d <= matchd3147d;
	-- d3149d
	sted3149d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3149d,
			Enable=>Enabled3149d,
			match=>matchd3149d,
			run=>run);

	reports(166) <= matchd3149d;
	Enabled3149d <= matchd3148d;
	-- d3150d
	sted3150d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3150d,
			Enable=>Enabled3150d,
			match=>matchd3150d,
			run=>run);

	-- d3151d
	sted3151d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3151d,
			Enable=>Enabled3151d,
			match=>matchd3151d,
			run=>run);

	Enabled3151d <= matchd3151d OR matchd3150d;
	-- d3152d
	sted3152d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3152d,
			Enable=>Enabled3152d,
			match=>matchd3152d,
			run=>run);

	Enabled3152d <= matchd3151d;
	-- d3153d
	sted3153d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3153d,
			Enable=>Enabled3153d,
			match=>matchd3153d,
			run=>run);

	Enabled3153d <= matchd3153d OR matchd3152d;
	-- d3154d
	sted3154d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3154d,
			Enable=>Enabled3154d,
			match=>matchd3154d,
			run=>run);

	Enabled3154d <= matchd3153d;
	-- d3155d
	sted3155d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3155d,
			Enable=>Enabled3155d,
			match=>matchd3155d,
			run=>run);

	Enabled3155d <= matchd3154d;
	-- d3156d
	sted3156d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3156d,
			Enable=>Enabled3156d,
			match=>matchd3156d,
			run=>run);

	Enabled3156d <= matchd3155d;
	-- d3157d
	sted3157d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3157d,
			Enable=>Enabled3157d,
			match=>matchd3157d,
			run=>run);

	Enabled3157d <= matchd3156d;
	-- d3158d
	sted3158d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3158d,
			Enable=>Enabled3158d,
			match=>matchd3158d,
			run=>run);

	Enabled3158d <= matchd3157d;
	-- d3159d
	sted3159d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3159d,
			Enable=>Enabled3159d,
			match=>matchd3159d,
			run=>run);

	Enabled3159d <= matchd3159d OR matchd3158d;
	-- d3160d
	sted3160d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3160d,
			Enable=>Enabled3160d,
			match=>matchd3160d,
			run=>run);

	Enabled3160d <= matchd3159d;
	-- d3161d
	sted3161d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3161d,
			Enable=>Enabled3161d,
			match=>matchd3161d,
			run=>run);

	Enabled3161d <= matchd3160d OR matchd3161d;
	-- d3162d
	sted3162d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3162d,
			Enable=>Enabled3162d,
			match=>matchd3162d,
			run=>run);

	Enabled3162d <= matchd3161d;
	-- d3163d
	sted3163d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3163d,
			Enable=>Enabled3163d,
			match=>matchd3163d,
			run=>run);

	Enabled3163d <= matchd3162d;
	-- d3164d
	sted3164d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3164d,
			Enable=>Enabled3164d,
			match=>matchd3164d,
			run=>run);

	Enabled3164d <= matchd3163d;
	-- d3165d
	sted3165d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3165d,
			Enable=>Enabled3165d,
			match=>matchd3165d,
			run=>run);

	Enabled3165d <= matchd3164d;
	-- d3166d
	sted3166d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3166d,
			Enable=>Enabled3166d,
			match=>matchd3166d,
			run=>run);

	-- d3167d
	sted3167d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3167d,
			Enable=>Enabled3167d,
			match=>matchd3167d,
			run=>run);

	Enabled3167d <= matchd3166d;
	-- d3168d
	sted3168d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3168d,
			Enable=>Enabled3168d,
			match=>matchd3168d,
			run=>run);

	Enabled3168d <= matchd3167d;
	-- d3169d
	sted3169d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3169d,
			Enable=>Enabled3169d,
			match=>matchd3169d,
			run=>run);

	Enabled3169d <= matchd3168d;
	-- d3170d
	sted3170d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3170d,
			Enable=>Enabled3170d,
			match=>matchd3170d,
			run=>run);

	Enabled3170d <= matchd3169d;
	-- d3171d
	sted3171d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3171d,
			Enable=>Enabled3171d,
			match=>matchd3171d,
			run=>run);

	Enabled3171d <= matchd3171d OR matchd3170d;
	-- d3172d
	sted3172d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3172d,
			Enable=>Enabled3172d,
			match=>matchd3172d,
			run=>run);

	Enabled3172d <= matchd3171d;
	-- d3173d
	sted3173d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3173d,
			Enable=>Enabled3173d,
			match=>matchd3173d,
			run=>run);

	Enabled3173d <= matchd3173d OR matchd3172d;
	-- d3174d
	sted3174d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3174d,
			Enable=>Enabled3174d,
			match=>matchd3174d,
			run=>run);

	Enabled3174d <= matchd3173d;
	-- d3175d
	sted3175d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3175d,
			Enable=>Enabled3175d,
			match=>matchd3175d,
			run=>run);

	Enabled3175d <= matchd3175d OR matchd3174d;
	-- d3176d
	sted3176d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3176d,
			Enable=>Enabled3176d,
			match=>matchd3176d,
			run=>run);

	Enabled3176d <= matchd3175d;
	-- d3177d
	sted3177d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3177d,
			Enable=>Enabled3177d,
			match=>matchd3177d,
			run=>run);

	Enabled3177d <= matchd3177d OR matchd3176d;
	-- d3178d
	sted3178d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3178d,
			Enable=>Enabled3178d,
			match=>matchd3178d,
			run=>run);

	Enabled3178d <= matchd3177d;
	-- d3179d
	sted3179d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3179d,
			Enable=>Enabled3179d,
			match=>matchd3179d,
			run=>run);

	Enabled3179d <= matchd3178d;
	-- d3180d
	sted3180d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3180d,
			Enable=>Enabled3180d,
			match=>matchd3180d,
			run=>run);

	Enabled3180d <= matchd3179d;
	-- d3181d
	sted3181d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3181d,
			Enable=>Enabled3181d,
			match=>matchd3181d,
			run=>run);

	Enabled3181d <= matchd3180d;
	-- d3183d
	sted3183d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3183d,
			Enable=>Enabled3183d,
			match=>matchd3183d,
			run=>run);

	-- d3184d
	sted3184d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3184d,
			Enable=>Enabled3184d,
			match=>matchd3184d,
			run=>run);

	Enabled3184d <= matchd3183d;
	-- d3185d
	sted3185d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3185d,
			Enable=>Enabled3185d,
			match=>matchd3185d,
			run=>run);

	Enabled3185d <= matchd3184d;
	-- d3186d
	sted3186d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3186d,
			Enable=>Enabled3186d,
			match=>matchd3186d,
			run=>run);

	Enabled3186d <= matchd3185d;
	-- d3187d
	sted3187d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3187d,
			Enable=>Enabled3187d,
			match=>matchd3187d,
			run=>run);

	Enabled3187d <= matchd3186d;
	-- d3188d
	sted3188d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3188d,
			Enable=>Enabled3188d,
			match=>matchd3188d,
			run=>run);

	Enabled3188d <= matchd3187d;
	-- d3189d
	sted3189d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3189d,
			Enable=>Enabled3189d,
			match=>matchd3189d,
			run=>run);

	Enabled3189d <= matchd3188d;
	-- d3190d
	sted3190d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3190d,
			Enable=>Enabled3190d,
			match=>matchd3190d,
			run=>run);

	Enabled3190d <= matchd3189d;
	-- d3191d
	sted3191d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3191d,
			Enable=>Enabled3191d,
			match=>matchd3191d,
			run=>run);

	Enabled3191d <= matchd3190d;
	-- d3192d
	sted3192d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3192d,
			Enable=>Enabled3192d,
			match=>matchd3192d,
			run=>run);

	Enabled3192d <= matchd3191d OR matchd3192d;
	-- d3193d
	sted3193d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3193d,
			Enable=>Enabled3193d,
			match=>matchd3193d,
			run=>run);

	Enabled3193d <= matchd3192d;
	-- d3194d
	sted3194d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3194d,
			Enable=>Enabled3194d,
			match=>matchd3194d,
			run=>run);

	Enabled3194d <= matchd3194d OR matchd3193d;
	-- d3195d
	sted3195d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3195d,
			Enable=>Enabled3195d,
			match=>matchd3195d,
			run=>run);

	Enabled3195d <= matchd3194d;
	-- d3196d
	sted3196d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3196d,
			Enable=>Enabled3196d,
			match=>matchd3196d,
			run=>run);

	Enabled3196d <= matchd3196d OR matchd3195d;
	-- d3197d
	sted3197d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3197d,
			Enable=>Enabled3197d,
			match=>matchd3197d,
			run=>run);

	Enabled3197d <= matchd3196d;
	-- d3198d
	sted3198d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3198d,
			Enable=>Enabled3198d,
			match=>matchd3198d,
			run=>run);

	Enabled3198d <= matchd3197d;
	-- d3199d
	sted3199d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3199d,
			Enable=>Enabled3199d,
			match=>matchd3199d,
			run=>run);

	Enabled3199d <= matchd3198d;
	-- d3200d
	sted3200d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3200d,
			Enable=>Enabled3200d,
			match=>matchd3200d,
			run=>run);

	Enabled3200d <= matchd3199d;
	-- d3201d
	sted3201d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3201d,
			Enable=>Enabled3201d,
			match=>matchd3201d,
			run=>run);

	reports(167) <= matchd3201d;
	Enabled3201d <= matchd3200d;
	-- d3202d
	sted3202d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3202d,
			Enable=>Enabled3202d,
			match=>matchd3202d,
			run=>run);

	-- d3203d
	sted3203d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3203d,
			Enable=>Enabled3203d,
			match=>matchd3203d,
			run=>run);

	Enabled3203d <= matchd3203d OR matchd3202d;
	-- d3204d
	sted3204d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3204d,
			Enable=>Enabled3204d,
			match=>matchd3204d,
			run=>run);

	Enabled3204d <= matchd3203d;
	-- d3205d
	sted3205d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3205d,
			Enable=>Enabled3205d,
			match=>matchd3205d,
			run=>run);

	Enabled3205d <= matchd3204d;
	-- d3206d
	sted3206d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3206d,
			Enable=>Enabled3206d,
			match=>matchd3206d,
			run=>run);

	Enabled3206d <= matchd3205d;
	-- d3207d
	sted3207d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3207d,
			Enable=>Enabled3207d,
			match=>matchd3207d,
			run=>run);

	Enabled3207d <= matchd3206d;
	-- d3208d
	sted3208d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3208d,
			Enable=>Enabled3208d,
			match=>matchd3208d,
			run=>run);

	Enabled3208d <= matchd3208d OR matchd3207d;
	-- d3209d
	sted3209d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3209d,
			Enable=>Enabled3209d,
			match=>matchd3209d,
			run=>run);

	Enabled3209d <= matchd3208d;
	-- d3210d
	sted3210d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3210d,
			Enable=>Enabled3210d,
			match=>matchd3210d,
			run=>run);

	Enabled3210d <= matchd3209d;
	-- d3211d
	sted3211d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3211d,
			Enable=>Enabled3211d,
			match=>matchd3211d,
			run=>run);

	Enabled3211d <= matchd3210d;
	-- d3212d
	sted3212d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3212d,
			Enable=>Enabled3212d,
			match=>matchd3212d,
			run=>run);

	Enabled3212d <= matchd3211d;
	-- d3213d
	sted3213d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3213d,
			Enable=>Enabled3213d,
			match=>matchd3213d,
			run=>run);

	reports(168) <= matchd3213d;
	Enabled3213d <= matchd3212d;
	-- d3214d
	sted3214d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3214d,
			Enable=>Enabled3214d,
			match=>matchd3214d,
			run=>run);

	-- d3215d
	sted3215d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3215d,
			Enable=>Enabled3215d,
			match=>matchd3215d,
			run=>run);

	Enabled3215d <= matchd3214d;
	-- d3216d
	sted3216d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3216d,
			Enable=>Enabled3216d,
			match=>matchd3216d,
			run=>run);

	Enabled3216d <= matchd3215d;
	-- d3217d
	sted3217d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3217d,
			Enable=>Enabled3217d,
			match=>matchd3217d,
			run=>run);

	Enabled3217d <= matchd3216d;
	-- d3218d
	sted3218d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3218d,
			Enable=>Enabled3218d,
			match=>matchd3218d,
			run=>run);

	Enabled3218d <= matchd3217d;
	-- d3219d
	sted3219d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3219d,
			Enable=>Enabled3219d,
			match=>matchd3219d,
			run=>run);

	Enabled3219d <= matchd3218d;
	-- d3220d
	sted3220d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3220d,
			Enable=>Enabled3220d,
			match=>matchd3220d,
			run=>run);

	Enabled3220d <= matchd3219d;
	-- d3221d
	sted3221d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3221d,
			Enable=>Enabled3221d,
			match=>matchd3221d,
			run=>run);

	Enabled3221d <= matchd3221d OR matchd3220d;
	-- d3222d
	sted3222d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3222d,
			Enable=>Enabled3222d,
			match=>matchd3222d,
			run=>run);

	Enabled3222d <= matchd3221d;
	-- d3223d
	sted3223d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3223d,
			Enable=>Enabled3223d,
			match=>matchd3223d,
			run=>run);

	Enabled3223d <= matchd3222d;
	-- d3224d
	sted3224d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3224d,
			Enable=>Enabled3224d,
			match=>matchd3224d,
			run=>run);

	Enabled3224d <= matchd3223d;
	-- d3225d
	sted3225d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3225d,
			Enable=>Enabled3225d,
			match=>matchd3225d,
			run=>run);

	Enabled3225d <= matchd3224d;
	-- d3226d
	sted3226d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3226d,
			Enable=>Enabled3226d,
			match=>matchd3226d,
			run=>run);

	reports(169) <= matchd3226d;
	Enabled3226d <= matchd3225d;
	-- d3227d
	sted3227d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3227d,
			Enable=>Enabled3227d,
			match=>matchd3227d,
			run=>run);

	-- d3228d
	sted3228d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3228d,
			Enable=>Enabled3228d,
			match=>matchd3228d,
			run=>run);

	Enabled3228d <= matchd3227d;
	-- d3229d
	sted3229d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3229d,
			Enable=>Enabled3229d,
			match=>matchd3229d,
			run=>run);

	Enabled3229d <= matchd3228d;
	-- d3230d
	sted3230d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3230d,
			Enable=>Enabled3230d,
			match=>matchd3230d,
			run=>run);

	Enabled3230d <= matchd3229d;
	-- d3231d
	sted3231d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3231d,
			Enable=>Enabled3231d,
			match=>matchd3231d,
			run=>run);

	Enabled3231d <= matchd3230d OR matchd3231d;
	-- d3232d
	sted3232d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3232d,
			Enable=>Enabled3232d,
			match=>matchd3232d,
			run=>run);

	Enabled3232d <= matchd3231d;
	-- d3233d
	sted3233d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3233d,
			Enable=>Enabled3233d,
			match=>matchd3233d,
			run=>run);

	Enabled3233d <= matchd3232d OR matchd3233d;
	-- d3234d
	sted3234d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3234d,
			Enable=>Enabled3234d,
			match=>matchd3234d,
			run=>run);

	Enabled3234d <= matchd3233d;
	-- d3235d
	sted3235d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3235d,
			Enable=>Enabled3235d,
			match=>matchd3235d,
			run=>run);

	Enabled3235d <= matchd3234d;
	-- d3236d
	sted3236d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3236d,
			Enable=>Enabled3236d,
			match=>matchd3236d,
			run=>run);

	Enabled3236d <= matchd3235d;
	-- d3237d
	sted3237d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3237d,
			Enable=>Enabled3237d,
			match=>matchd3237d,
			run=>run);

	reports(170) <= matchd3237d;
	Enabled3237d <= matchd3236d;
	-- d3238d
	sted3238d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3238d,
			Enable=>Enabled3238d,
			match=>matchd3238d,
			run=>run);

	-- d3239d
	sted3239d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3239d,
			Enable=>Enabled3239d,
			match=>matchd3239d,
			run=>run);

	Enabled3239d <= matchd3238d;
	-- d3240d
	sted3240d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3240d,
			Enable=>Enabled3240d,
			match=>matchd3240d,
			run=>run);

	Enabled3240d <= matchd3239d;
	-- d3241d
	sted3241d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3241d,
			Enable=>Enabled3241d,
			match=>matchd3241d,
			run=>run);

	Enabled3241d <= matchd3240d;
	-- d3242d
	sted3242d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3242d,
			Enable=>Enabled3242d,
			match=>matchd3242d,
			run=>run);

	Enabled3242d <= matchd3241d;
	-- d3243d
	sted3243d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3243d,
			Enable=>Enabled3243d,
			match=>matchd3243d,
			run=>run);

	Enabled3243d <= matchd3242d;
	-- d3244d
	sted3244d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3244d,
			Enable=>Enabled3244d,
			match=>matchd3244d,
			run=>run);

	reports(171) <= matchd3244d;
	Enabled3244d <= matchd3243d;
	-- d3245d
	sted3245d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3245d,
			Enable=>Enabled3245d,
			match=>matchd3245d,
			run=>run);

	-- d3246d
	sted3246d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3246d,
			Enable=>Enabled3246d,
			match=>matchd3246d,
			run=>run);

	Enabled3246d <= matchd3246d OR matchd3245d;
	-- d3247d
	sted3247d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3247d,
			Enable=>Enabled3247d,
			match=>matchd3247d,
			run=>run);

	Enabled3247d <= matchd3246d;
	-- d3248d
	sted3248d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3248d,
			Enable=>Enabled3248d,
			match=>matchd3248d,
			run=>run);

	Enabled3248d <= matchd3247d;
	-- d3249d
	sted3249d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3249d,
			Enable=>Enabled3249d,
			match=>matchd3249d,
			run=>run);

	Enabled3249d <= matchd3248d;
	-- d3250d
	sted3250d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3250d,
			Enable=>Enabled3250d,
			match=>matchd3250d,
			run=>run);

	Enabled3250d <= matchd3249d;
	-- d3251d
	sted3251d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3251d,
			Enable=>Enabled3251d,
			match=>matchd3251d,
			run=>run);

	Enabled3251d <= matchd3250d OR matchd3251d;
	-- d3252d
	sted3252d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3252d,
			Enable=>Enabled3252d,
			match=>matchd3252d,
			run=>run);

	Enabled3252d <= matchd3251d;
	-- d3253d
	sted3253d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3253d,
			Enable=>Enabled3253d,
			match=>matchd3253d,
			run=>run);

	Enabled3253d <= matchd3252d;
	-- d3254d
	sted3254d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3254d,
			Enable=>Enabled3254d,
			match=>matchd3254d,
			run=>run);

	Enabled3254d <= matchd3253d;
	-- d3255d
	sted3255d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3255d,
			Enable=>Enabled3255d,
			match=>matchd3255d,
			run=>run);

	Enabled3255d <= matchd3254d;
	-- d3256d
	sted3256d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3256d,
			Enable=>Enabled3256d,
			match=>matchd3256d,
			run=>run);

	Enabled3256d <= matchd3255d;
	-- d3257d
	sted3257d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3257d,
			Enable=>Enabled3257d,
			match=>matchd3257d,
			run=>run);

	Enabled3257d <= matchd3256d OR matchd3257d;
	-- d3258d
	sted3258d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3258d,
			Enable=>Enabled3258d,
			match=>matchd3258d,
			run=>run);

	Enabled3258d <= matchd3257d;
	-- d3259d
	sted3259d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3259d,
			Enable=>Enabled3259d,
			match=>matchd3259d,
			run=>run);

	Enabled3259d <= matchd3258d;
	-- d3260d
	sted3260d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3260d,
			Enable=>Enabled3260d,
			match=>matchd3260d,
			run=>run);

	reports(172) <= matchd3260d;
	Enabled3260d <= matchd3259d;
	-- d3261d
	sted3261d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3261d,
			Enable=>Enabled3261d,
			match=>matchd3261d,
			run=>run);

	-- d3262d
	sted3262d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3262d,
			Enable=>Enabled3262d,
			match=>matchd3262d,
			run=>run);

	Enabled3262d <= matchd3261d OR matchd3262d;
	-- d3263d
	sted3263d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3263d,
			Enable=>Enabled3263d,
			match=>matchd3263d,
			run=>run);

	Enabled3263d <= matchd3262d;
	-- d3264d
	sted3264d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3264d,
			Enable=>Enabled3264d,
			match=>matchd3264d,
			run=>run);

	Enabled3264d <= matchd3263d OR matchd3264d;
	-- d3265d
	sted3265d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3265d,
			Enable=>Enabled3265d,
			match=>matchd3265d,
			run=>run);

	Enabled3265d <= matchd3264d;
	-- d3266d
	sted3266d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3266d,
			Enable=>Enabled3266d,
			match=>matchd3266d,
			run=>run);

	Enabled3266d <= matchd3265d;
	-- d3267d
	sted3267d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3267d,
			Enable=>Enabled3267d,
			match=>matchd3267d,
			run=>run);

	Enabled3267d <= matchd3266d;
	-- d3268d
	sted3268d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3268d,
			Enable=>Enabled3268d,
			match=>matchd3268d,
			run=>run);

	Enabled3268d <= matchd3267d;
	-- d3269d
	sted3269d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3269d,
			Enable=>Enabled3269d,
			match=>matchd3269d,
			run=>run);

	Enabled3269d <= matchd3268d;
	-- d3270d
	sted3270d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3270d,
			Enable=>Enabled3270d,
			match=>matchd3270d,
			run=>run);

	Enabled3270d <= matchd3270d OR matchd3269d;
	-- d3271d
	sted3271d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3271d,
			Enable=>Enabled3271d,
			match=>matchd3271d,
			run=>run);

	Enabled3271d <= matchd3270d;
	-- d3272d
	sted3272d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3272d,
			Enable=>Enabled3272d,
			match=>matchd3272d,
			run=>run);

	Enabled3272d <= matchd3272d OR matchd3271d;
	-- d3273d
	sted3273d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3273d,
			Enable=>Enabled3273d,
			match=>matchd3273d,
			run=>run);

	Enabled3273d <= matchd3272d;
	-- d3274d
	sted3274d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3274d,
			Enable=>Enabled3274d,
			match=>matchd3274d,
			run=>run);

	Enabled3274d <= matchd3273d;
	-- d3275d
	sted3275d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3275d,
			Enable=>Enabled3275d,
			match=>matchd3275d,
			run=>run);

	Enabled3275d <= matchd3274d;
	-- d3276d
	sted3276d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3276d,
			Enable=>Enabled3276d,
			match=>matchd3276d,
			run=>run);

	Enabled3276d <= matchd3275d;
	-- d3277d
	sted3277d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3277d,
			Enable=>Enabled3277d,
			match=>matchd3277d,
			run=>run);

	Enabled3277d <= matchd3276d;
	-- d3278d
	sted3278d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3278d,
			Enable=>Enabled3278d,
			match=>matchd3278d,
			run=>run);

	-- d3279d
	sted3279d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3279d,
			Enable=>Enabled3279d,
			match=>matchd3279d,
			run=>run);

	Enabled3279d <= matchd3278d;
	-- d3280d
	sted3280d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3280d,
			Enable=>Enabled3280d,
			match=>matchd3280d,
			run=>run);

	Enabled3280d <= matchd3279d;
	-- d3281d
	sted3281d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3281d,
			Enable=>Enabled3281d,
			match=>matchd3281d,
			run=>run);

	Enabled3281d <= matchd3280d;
	-- d3282d
	sted3282d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3282d,
			Enable=>Enabled3282d,
			match=>matchd3282d,
			run=>run);

	Enabled3282d <= matchd3281d;
	-- d3283d
	sted3283d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3283d,
			Enable=>Enabled3283d,
			match=>matchd3283d,
			run=>run);

	Enabled3283d <= matchd3283d OR matchd3282d;
	-- d3284d
	sted3284d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3284d,
			Enable=>Enabled3284d,
			match=>matchd3284d,
			run=>run);

	Enabled3284d <= matchd3283d;
	-- d3285d
	sted3285d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3285d,
			Enable=>Enabled3285d,
			match=>matchd3285d,
			run=>run);

	Enabled3285d <= matchd3285d OR matchd3284d;
	-- d3286d
	sted3286d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3286d,
			Enable=>Enabled3286d,
			match=>matchd3286d,
			run=>run);

	Enabled3286d <= matchd3285d;
	-- d3287d
	sted3287d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3287d,
			Enable=>Enabled3287d,
			match=>matchd3287d,
			run=>run);

	Enabled3287d <= matchd3286d OR matchd3287d;
	-- d3288d
	sted3288d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3288d,
			Enable=>Enabled3288d,
			match=>matchd3288d,
			run=>run);

	Enabled3288d <= matchd3287d;
	-- d3289d
	sted3289d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3289d,
			Enable=>Enabled3289d,
			match=>matchd3289d,
			run=>run);

	Enabled3289d <= matchd3289d OR matchd3288d;
	-- d3290d
	sted3290d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3290d,
			Enable=>Enabled3290d,
			match=>matchd3290d,
			run=>run);

	Enabled3290d <= matchd3289d;
	-- d3291d
	sted3291d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3291d,
			Enable=>Enabled3291d,
			match=>matchd3291d,
			run=>run);

	Enabled3291d <= matchd3290d;
	-- d3292d
	sted3292d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3292d,
			Enable=>Enabled3292d,
			match=>matchd3292d,
			run=>run);

	Enabled3292d <= matchd3291d;
	-- d3293d
	sted3293d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3293d,
			Enable=>Enabled3293d,
			match=>matchd3293d,
			run=>run);

	Enabled3293d <= matchd3292d;
	-- d3294d
	sted3294d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3294d,
			Enable=>Enabled3294d,
			match=>matchd3294d,
			run=>run);

	Enabled3294d <= matchd3293d;
	-- d3296d
	sted3296d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3296d,
			Enable=>Enabled3296d,
			match=>matchd3296d,
			run=>run);

	-- d3297d
	sted3297d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3297d,
			Enable=>Enabled3297d,
			match=>matchd3297d,
			run=>run);

	Enabled3297d <= matchd3296d;
	-- d3298d
	sted3298d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3298d,
			Enable=>Enabled3298d,
			match=>matchd3298d,
			run=>run);

	Enabled3298d <= matchd3297d;
	-- d3299d
	sted3299d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3299d,
			Enable=>Enabled3299d,
			match=>matchd3299d,
			run=>run);

	Enabled3299d <= matchd3298d;
	-- d3300d
	sted3300d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3300d,
			Enable=>Enabled3300d,
			match=>matchd3300d,
			run=>run);

	Enabled3300d <= matchd3299d;
	-- d3301d
	sted3301d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3301d,
			Enable=>Enabled3301d,
			match=>matchd3301d,
			run=>run);

	Enabled3301d <= matchd3300d;
	-- d3302d
	sted3302d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3302d,
			Enable=>Enabled3302d,
			match=>matchd3302d,
			run=>run);

	Enabled3302d <= matchd3301d OR matchd3302d;
	-- d3303d
	sted3303d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3303d,
			Enable=>Enabled3303d,
			match=>matchd3303d,
			run=>run);

	Enabled3303d <= matchd3302d;
	-- d3304d
	sted3304d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3304d,
			Enable=>Enabled3304d,
			match=>matchd3304d,
			run=>run);

	Enabled3304d <= matchd3304d OR matchd3303d;
	-- d3305d
	sted3305d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3305d,
			Enable=>Enabled3305d,
			match=>matchd3305d,
			run=>run);

	Enabled3305d <= matchd3304d;
	-- d3306d
	sted3306d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3306d,
			Enable=>Enabled3306d,
			match=>matchd3306d,
			run=>run);

	Enabled3306d <= matchd3305d;
	-- d3307d
	sted3307d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3307d,
			Enable=>Enabled3307d,
			match=>matchd3307d,
			run=>run);

	Enabled3307d <= matchd3306d;
	-- d3308d
	sted3308d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3308d,
			Enable=>Enabled3308d,
			match=>matchd3308d,
			run=>run);

	Enabled3308d <= matchd3307d;
	-- d3309d
	sted3309d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3309d,
			Enable=>Enabled3309d,
			match=>matchd3309d,
			run=>run);

	reports(173) <= matchd3309d;
	Enabled3309d <= matchd3308d;
	-- d3310d
	sted3310d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3310d,
			Enable=>Enabled3310d,
			match=>matchd3310d,
			run=>run);

	-- d3311d
	sted3311d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3311d,
			Enable=>Enabled3311d,
			match=>matchd3311d,
			run=>run);

	Enabled3311d <= matchd3310d OR matchd3311d;
	-- d3312d
	sted3312d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3312d,
			Enable=>Enabled3312d,
			match=>matchd3312d,
			run=>run);

	Enabled3312d <= matchd3311d;
	-- d3313d
	sted3313d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3313d,
			Enable=>Enabled3313d,
			match=>matchd3313d,
			run=>run);

	Enabled3313d <= matchd3312d;
	-- d3314d
	sted3314d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3314d,
			Enable=>Enabled3314d,
			match=>matchd3314d,
			run=>run);

	Enabled3314d <= matchd3313d;
	-- d3315d
	sted3315d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3315d,
			Enable=>Enabled3315d,
			match=>matchd3315d,
			run=>run);

	Enabled3315d <= matchd3314d;
	-- d3316d
	sted3316d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3316d,
			Enable=>Enabled3316d,
			match=>matchd3316d,
			run=>run);

	Enabled3316d <= matchd3315d;
	-- d3317d
	sted3317d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3317d,
			Enable=>Enabled3317d,
			match=>matchd3317d,
			run=>run);

	Enabled3317d <= matchd3316d;
	-- d3318d
	sted3318d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3318d,
			Enable=>Enabled3318d,
			match=>matchd3318d,
			run=>run);

	Enabled3318d <= matchd3317d;
	-- d3319d
	sted3319d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3319d,
			Enable=>Enabled3319d,
			match=>matchd3319d,
			run=>run);

	Enabled3319d <= matchd3318d;
	-- d3320d
	sted3320d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3320d,
			Enable=>Enabled3320d,
			match=>matchd3320d,
			run=>run);

	Enabled3320d <= matchd3319d;
	-- d3321d
	sted3321d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3321d,
			Enable=>Enabled3321d,
			match=>matchd3321d,
			run=>run);

	Enabled3321d <= matchd3320d;
	-- d3322d
	sted3322d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3322d,
			Enable=>Enabled3322d,
			match=>matchd3322d,
			run=>run);

	Enabled3322d <= matchd3321d;
	-- d3323d
	sted3323d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3323d,
			Enable=>Enabled3323d,
			match=>matchd3323d,
			run=>run);

	reports(174) <= matchd3323d;
	Enabled3323d <= matchd3322d;
	-- d3324d
	sted3324d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3324d,
			Enable=>Enabled3324d,
			match=>matchd3324d,
			run=>run);

	-- d3325d
	sted3325d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3325d,
			Enable=>Enabled3325d,
			match=>matchd3325d,
			run=>run);

	Enabled3325d <= matchd3324d OR matchd3325d;
	-- d3326d
	sted3326d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3326d,
			Enable=>Enabled3326d,
			match=>matchd3326d,
			run=>run);

	Enabled3326d <= matchd3325d;
	-- d3327d
	sted3327d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3327d,
			Enable=>Enabled3327d,
			match=>matchd3327d,
			run=>run);

	Enabled3327d <= matchd3326d;
	-- d3328d
	sted3328d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3328d,
			Enable=>Enabled3328d,
			match=>matchd3328d,
			run=>run);

	Enabled3328d <= matchd3327d;
	-- d3329d
	sted3329d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3329d,
			Enable=>Enabled3329d,
			match=>matchd3329d,
			run=>run);

	Enabled3329d <= matchd3328d;
	-- d3330d
	sted3330d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3330d,
			Enable=>Enabled3330d,
			match=>matchd3330d,
			run=>run);

	Enabled3330d <= matchd3329d OR matchd3330d;
	-- d3331d
	sted3331d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3331d,
			Enable=>Enabled3331d,
			match=>matchd3331d,
			run=>run);

	Enabled3331d <= matchd3330d;
	-- d3332d
	sted3332d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3332d,
			Enable=>Enabled3332d,
			match=>matchd3332d,
			run=>run);

	Enabled3332d <= matchd3331d;
	-- d3333d
	sted3333d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3333d,
			Enable=>Enabled3333d,
			match=>matchd3333d,
			run=>run);

	Enabled3333d <= matchd3332d;
	-- d3334d
	sted3334d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3334d,
			Enable=>Enabled3334d,
			match=>matchd3334d,
			run=>run);

	reports(175) <= matchd3334d;
	Enabled3334d <= matchd3333d;
	-- d3335d
	sted3335d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3335d,
			Enable=>Enabled3335d,
			match=>matchd3335d,
			run=>run);

	-- d3336d
	sted3336d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3336d,
			Enable=>Enabled3336d,
			match=>matchd3336d,
			run=>run);

	Enabled3336d <= matchd3336d OR matchd3335d;
	-- d3337d
	sted3337d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3337d,
			Enable=>Enabled3337d,
			match=>matchd3337d,
			run=>run);

	Enabled3337d <= matchd3336d;
	-- d3338d
	sted3338d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3338d,
			Enable=>Enabled3338d,
			match=>matchd3338d,
			run=>run);

	Enabled3338d <= matchd3337d;
	-- d3339d
	sted3339d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3339d,
			Enable=>Enabled3339d,
			match=>matchd3339d,
			run=>run);

	Enabled3339d <= matchd3338d;
	-- d3340d
	sted3340d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3340d,
			Enable=>Enabled3340d,
			match=>matchd3340d,
			run=>run);

	Enabled3340d <= matchd3339d;
	-- d3341d
	sted3341d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3341d,
			Enable=>Enabled3341d,
			match=>matchd3341d,
			run=>run);

	Enabled3341d <= matchd3340d;
	-- d3342d
	sted3342d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3342d,
			Enable=>Enabled3342d,
			match=>matchd3342d,
			run=>run);

	Enabled3342d <= matchd3342d OR matchd3341d;
	-- d3343d
	sted3343d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3343d,
			Enable=>Enabled3343d,
			match=>matchd3343d,
			run=>run);

	Enabled3343d <= matchd3342d;
	-- d3344d
	sted3344d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3344d,
			Enable=>Enabled3344d,
			match=>matchd3344d,
			run=>run);

	Enabled3344d <= matchd3343d;
	-- d3345d
	sted3345d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3345d,
			Enable=>Enabled3345d,
			match=>matchd3345d,
			run=>run);

	Enabled3345d <= matchd3344d;
	-- d3346d
	sted3346d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3346d,
			Enable=>Enabled3346d,
			match=>matchd3346d,
			run=>run);

	Enabled3346d <= matchd3345d;
	-- d3347d
	sted3347d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3347d,
			Enable=>Enabled3347d,
			match=>matchd3347d,
			run=>run);

	reports(176) <= matchd3347d;
	Enabled3347d <= matchd3346d;
	-- d3348d
	sted3348d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3348d,
			Enable=>Enabled3348d,
			match=>matchd3348d,
			run=>run);

	-- d3349d
	sted3349d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3349d,
			Enable=>Enabled3349d,
			match=>matchd3349d,
			run=>run);

	Enabled3349d <= matchd3348d OR matchd3349d;
	-- d3350d
	sted3350d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3350d,
			Enable=>Enabled3350d,
			match=>matchd3350d,
			run=>run);

	Enabled3350d <= matchd3349d;
	-- d3351d
	sted3351d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3351d,
			Enable=>Enabled3351d,
			match=>matchd3351d,
			run=>run);

	Enabled3351d <= matchd3350d;
	-- d3352d
	sted3352d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3352d,
			Enable=>Enabled3352d,
			match=>matchd3352d,
			run=>run);

	Enabled3352d <= matchd3351d;
	-- d3353d
	sted3353d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3353d,
			Enable=>Enabled3353d,
			match=>matchd3353d,
			run=>run);

	Enabled3353d <= matchd3352d;
	-- d3354d
	sted3354d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3354d,
			Enable=>Enabled3354d,
			match=>matchd3354d,
			run=>run);

	Enabled3354d <= matchd3353d;
	-- d3355d
	sted3355d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3355d,
			Enable=>Enabled3355d,
			match=>matchd3355d,
			run=>run);

	Enabled3355d <= matchd3354d;
	-- d3356d
	sted3356d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3356d,
			Enable=>Enabled3356d,
			match=>matchd3356d,
			run=>run);

	Enabled3356d <= matchd3355d OR matchd3356d;
	-- d3357d
	sted3357d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3357d,
			Enable=>Enabled3357d,
			match=>matchd3357d,
			run=>run);

	Enabled3357d <= matchd3356d;
	-- d3358d
	sted3358d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3358d,
			Enable=>Enabled3358d,
			match=>matchd3358d,
			run=>run);

	Enabled3358d <= matchd3357d;
	-- d3359d
	sted3359d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3359d,
			Enable=>Enabled3359d,
			match=>matchd3359d,
			run=>run);

	Enabled3359d <= matchd3358d;
	-- d3360d
	sted3360d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3360d,
			Enable=>Enabled3360d,
			match=>matchd3360d,
			run=>run);

	Enabled3360d <= matchd3359d;
	-- d3361d
	sted3361d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3361d,
			Enable=>Enabled3361d,
			match=>matchd3361d,
			run=>run);

	reports(177) <= matchd3361d;
	Enabled3361d <= matchd3360d;
	-- d3362d
	sted3362d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3362d,
			Enable=>Enabled3362d,
			match=>matchd3362d,
			run=>run);

	-- d3363d
	sted3363d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3363d,
			Enable=>Enabled3363d,
			match=>matchd3363d,
			run=>run);

	Enabled3363d <= matchd3363d OR matchd3362d;
	-- d3364d
	sted3364d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3364d,
			Enable=>Enabled3364d,
			match=>matchd3364d,
			run=>run);

	Enabled3364d <= matchd3363d;
	-- d3365d
	sted3365d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3365d,
			Enable=>Enabled3365d,
			match=>matchd3365d,
			run=>run);

	Enabled3365d <= matchd3364d;
	-- d3366d
	sted3366d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3366d,
			Enable=>Enabled3366d,
			match=>matchd3366d,
			run=>run);

	Enabled3366d <= matchd3365d;
	-- d3367d
	sted3367d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3367d,
			Enable=>Enabled3367d,
			match=>matchd3367d,
			run=>run);

	Enabled3367d <= matchd3366d;
	-- d3368d
	sted3368d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3368d,
			Enable=>Enabled3368d,
			match=>matchd3368d,
			run=>run);

	Enabled3368d <= matchd3367d OR matchd3368d;
	-- d3369d
	sted3369d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3369d,
			Enable=>Enabled3369d,
			match=>matchd3369d,
			run=>run);

	Enabled3369d <= matchd3368d;
	-- d3370d
	sted3370d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3370d,
			Enable=>Enabled3370d,
			match=>matchd3370d,
			run=>run);

	Enabled3370d <= matchd3369d;
	-- d3371d
	sted3371d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3371d,
			Enable=>Enabled3371d,
			match=>matchd3371d,
			run=>run);

	Enabled3371d <= matchd3370d;
	-- d3372d
	sted3372d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3372d,
			Enable=>Enabled3372d,
			match=>matchd3372d,
			run=>run);

	Enabled3372d <= matchd3371d;
	-- d3373d
	sted3373d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3373d,
			Enable=>Enabled3373d,
			match=>matchd3373d,
			run=>run);

	Enabled3373d <= matchd3372d OR matchd3373d;
	-- d3374d
	sted3374d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3374d,
			Enable=>Enabled3374d,
			match=>matchd3374d,
			run=>run);

	Enabled3374d <= matchd3373d;
	-- d3375d
	sted3375d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3375d,
			Enable=>Enabled3375d,
			match=>matchd3375d,
			run=>run);

	Enabled3375d <= matchd3374d;
	-- d3376d
	sted3376d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3376d,
			Enable=>Enabled3376d,
			match=>matchd3376d,
			run=>run);

	Enabled3376d <= matchd3375d;
	-- d3377d
	sted3377d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3377d,
			Enable=>Enabled3377d,
			match=>matchd3377d,
			run=>run);

	reports(178) <= matchd3377d;
	Enabled3377d <= matchd3376d;
	-- d3378d
	sted3378d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3378d,
			Enable=>Enabled3378d,
			match=>matchd3378d,
			run=>run);

	-- d3379d
	sted3379d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3379d,
			Enable=>Enabled3379d,
			match=>matchd3379d,
			run=>run);

	Enabled3379d <= matchd3378d OR matchd3379d;
	-- d3380d
	sted3380d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3380d,
			Enable=>Enabled3380d,
			match=>matchd3380d,
			run=>run);

	Enabled3380d <= matchd3379d;
	-- d3381d
	sted3381d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3381d,
			Enable=>Enabled3381d,
			match=>matchd3381d,
			run=>run);

	Enabled3381d <= matchd3380d;
	-- d3382d
	sted3382d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3382d,
			Enable=>Enabled3382d,
			match=>matchd3382d,
			run=>run);

	Enabled3382d <= matchd3381d;
	-- d3383d
	sted3383d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3383d,
			Enable=>Enabled3383d,
			match=>matchd3383d,
			run=>run);

	Enabled3383d <= matchd3382d;
	-- d3384d
	sted3384d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3384d,
			Enable=>Enabled3384d,
			match=>matchd3384d,
			run=>run);

	Enabled3384d <= matchd3384d OR matchd3383d;
	-- d3385d
	sted3385d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3385d,
			Enable=>Enabled3385d,
			match=>matchd3385d,
			run=>run);

	Enabled3385d <= matchd3384d;
	-- d3386d
	sted3386d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3386d,
			Enable=>Enabled3386d,
			match=>matchd3386d,
			run=>run);

	Enabled3386d <= matchd3385d;
	-- d3387d
	sted3387d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3387d,
			Enable=>Enabled3387d,
			match=>matchd3387d,
			run=>run);

	Enabled3387d <= matchd3386d;
	-- d3388d
	sted3388d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3388d,
			Enable=>Enabled3388d,
			match=>matchd3388d,
			run=>run);

	reports(179) <= matchd3388d;
	Enabled3388d <= matchd3387d;
	-- d3389d
	sted3389d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3389d,
			Enable=>Enabled3389d,
			match=>matchd3389d,
			run=>run);

	-- d3390d
	sted3390d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3390d,
			Enable=>Enabled3390d,
			match=>matchd3390d,
			run=>run);

	Enabled3390d <= matchd3389d OR matchd3390d;
	-- d3391d
	sted3391d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3391d,
			Enable=>Enabled3391d,
			match=>matchd3391d,
			run=>run);

	Enabled3391d <= matchd3390d;
	-- d3392d
	sted3392d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3392d,
			Enable=>Enabled3392d,
			match=>matchd3392d,
			run=>run);

	Enabled3392d <= matchd3391d;
	-- d3393d
	sted3393d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3393d,
			Enable=>Enabled3393d,
			match=>matchd3393d,
			run=>run);

	Enabled3393d <= matchd3392d;
	-- d3394d
	sted3394d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3394d,
			Enable=>Enabled3394d,
			match=>matchd3394d,
			run=>run);

	Enabled3394d <= matchd3393d;
	-- d3395d
	sted3395d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3395d,
			Enable=>Enabled3395d,
			match=>matchd3395d,
			run=>run);

	Enabled3395d <= matchd3395d OR matchd3394d;
	-- d3396d
	sted3396d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3396d,
			Enable=>Enabled3396d,
			match=>matchd3396d,
			run=>run);

	Enabled3396d <= matchd3395d;
	-- d3397d
	sted3397d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3397d,
			Enable=>Enabled3397d,
			match=>matchd3397d,
			run=>run);

	Enabled3397d <= matchd3396d;
	-- d3398d
	sted3398d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3398d,
			Enable=>Enabled3398d,
			match=>matchd3398d,
			run=>run);

	Enabled3398d <= matchd3397d;
	-- d3399d
	sted3399d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3399d,
			Enable=>Enabled3399d,
			match=>matchd3399d,
			run=>run);

	reports(180) <= matchd3399d;
	Enabled3399d <= matchd3398d;
	-- d3400d
	sted3400d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3400d,
			Enable=>Enabled3400d,
			match=>matchd3400d,
			run=>run);

	-- d3401d
	sted3401d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3401d,
			Enable=>Enabled3401d,
			match=>matchd3401d,
			run=>run);

	Enabled3401d <= matchd3401d OR matchd3400d;
	-- d3402d
	sted3402d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3402d,
			Enable=>Enabled3402d,
			match=>matchd3402d,
			run=>run);

	Enabled3402d <= matchd3401d;
	-- d3403d
	sted3403d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3403d,
			Enable=>Enabled3403d,
			match=>matchd3403d,
			run=>run);

	Enabled3403d <= matchd3402d;
	-- d3404d
	sted3404d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3404d,
			Enable=>Enabled3404d,
			match=>matchd3404d,
			run=>run);

	Enabled3404d <= matchd3403d;
	-- d3405d
	sted3405d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3405d,
			Enable=>Enabled3405d,
			match=>matchd3405d,
			run=>run);

	Enabled3405d <= matchd3404d;
	-- d3406d
	sted3406d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3406d,
			Enable=>Enabled3406d,
			match=>matchd3406d,
			run=>run);

	Enabled3406d <= matchd3405d OR matchd3406d;
	-- d3407d
	sted3407d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3407d,
			Enable=>Enabled3407d,
			match=>matchd3407d,
			run=>run);

	Enabled3407d <= matchd3406d;
	-- d3408d
	sted3408d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3408d,
			Enable=>Enabled3408d,
			match=>matchd3408d,
			run=>run);

	Enabled3408d <= matchd3407d;
	-- d3409d
	sted3409d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3409d,
			Enable=>Enabled3409d,
			match=>matchd3409d,
			run=>run);

	Enabled3409d <= matchd3408d;
	-- d3410d
	sted3410d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3410d,
			Enable=>Enabled3410d,
			match=>matchd3410d,
			run=>run);

	Enabled3410d <= matchd3409d;
	-- d3411d
	sted3411d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3411d,
			Enable=>Enabled3411d,
			match=>matchd3411d,
			run=>run);

	reports(181) <= matchd3411d;
	Enabled3411d <= matchd3410d;
	-- d3412d
	sted3412d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3412d,
			Enable=>Enabled3412d,
			match=>matchd3412d,
			run=>run);

	-- d3413d
	sted3413d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3413d,
			Enable=>Enabled3413d,
			match=>matchd3413d,
			run=>run);

	Enabled3413d <= matchd3412d OR matchd3413d;
	-- d3414d
	sted3414d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3414d,
			Enable=>Enabled3414d,
			match=>matchd3414d,
			run=>run);

	Enabled3414d <= matchd3413d;
	-- d3415d
	sted3415d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3415d,
			Enable=>Enabled3415d,
			match=>matchd3415d,
			run=>run);

	Enabled3415d <= matchd3414d;
	-- d3416d
	sted3416d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3416d,
			Enable=>Enabled3416d,
			match=>matchd3416d,
			run=>run);

	Enabled3416d <= matchd3415d;
	-- d3417d
	sted3417d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3417d,
			Enable=>Enabled3417d,
			match=>matchd3417d,
			run=>run);

	Enabled3417d <= matchd3416d;
	-- d3418d
	sted3418d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3418d,
			Enable=>Enabled3418d,
			match=>matchd3418d,
			run=>run);

	Enabled3418d <= matchd3417d;
	-- d3419d
	sted3419d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3419d,
			Enable=>Enabled3419d,
			match=>matchd3419d,
			run=>run);

	Enabled3419d <= matchd3419d OR matchd3418d;
	-- d3420d
	sted3420d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3420d,
			Enable=>Enabled3420d,
			match=>matchd3420d,
			run=>run);

	Enabled3420d <= matchd3419d;
	-- d3421d
	sted3421d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3421d,
			Enable=>Enabled3421d,
			match=>matchd3421d,
			run=>run);

	Enabled3421d <= matchd3420d;
	-- d3422d
	sted3422d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3422d,
			Enable=>Enabled3422d,
			match=>matchd3422d,
			run=>run);

	Enabled3422d <= matchd3421d;
	-- d3423d
	sted3423d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3423d,
			Enable=>Enabled3423d,
			match=>matchd3423d,
			run=>run);

	reports(182) <= matchd3423d;
	Enabled3423d <= matchd3422d;
	-- d3424d
	sted3424d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3424d,
			Enable=>Enabled3424d,
			match=>matchd3424d,
			run=>run);

	-- d3425d
	sted3425d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3425d,
			Enable=>Enabled3425d,
			match=>matchd3425d,
			run=>run);

	Enabled3425d <= matchd3425d OR matchd3424d;
	-- d3426d
	sted3426d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3426d,
			Enable=>Enabled3426d,
			match=>matchd3426d,
			run=>run);

	Enabled3426d <= matchd3425d;
	-- d3427d
	sted3427d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3427d,
			Enable=>Enabled3427d,
			match=>matchd3427d,
			run=>run);

	Enabled3427d <= matchd3426d;
	-- d3428d
	sted3428d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3428d,
			Enable=>Enabled3428d,
			match=>matchd3428d,
			run=>run);

	Enabled3428d <= matchd3427d;
	-- d3429d
	sted3429d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3429d,
			Enable=>Enabled3429d,
			match=>matchd3429d,
			run=>run);

	Enabled3429d <= matchd3428d;
	-- d3430d
	sted3430d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3430d,
			Enable=>Enabled3430d,
			match=>matchd3430d,
			run=>run);

	Enabled3430d <= matchd3429d OR matchd3430d;
	-- d3431d
	sted3431d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3431d,
			Enable=>Enabled3431d,
			match=>matchd3431d,
			run=>run);

	Enabled3431d <= matchd3430d;
	-- d3432d
	sted3432d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3432d,
			Enable=>Enabled3432d,
			match=>matchd3432d,
			run=>run);

	Enabled3432d <= matchd3431d;
	-- d3433d
	sted3433d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3433d,
			Enable=>Enabled3433d,
			match=>matchd3433d,
			run=>run);

	Enabled3433d <= matchd3432d;
	-- d3434d
	sted3434d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3434d,
			Enable=>Enabled3434d,
			match=>matchd3434d,
			run=>run);

	Enabled3434d <= matchd3433d;
	-- d3435d
	sted3435d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3435d,
			Enable=>Enabled3435d,
			match=>matchd3435d,
			run=>run);

	reports(183) <= matchd3435d;
	Enabled3435d <= matchd3434d;
	-- d3436d
	sted3436d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3436d,
			Enable=>Enabled3436d,
			match=>matchd3436d,
			run=>run);

	-- d3437d
	sted3437d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3437d,
			Enable=>Enabled3437d,
			match=>matchd3437d,
			run=>run);

	Enabled3437d <= matchd3436d OR matchd3437d;
	-- d3438d
	sted3438d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3438d,
			Enable=>Enabled3438d,
			match=>matchd3438d,
			run=>run);

	Enabled3438d <= matchd3437d;
	-- d3439d
	sted3439d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3439d,
			Enable=>Enabled3439d,
			match=>matchd3439d,
			run=>run);

	Enabled3439d <= matchd3438d;
	-- d3440d
	sted3440d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3440d,
			Enable=>Enabled3440d,
			match=>matchd3440d,
			run=>run);

	Enabled3440d <= matchd3439d;
	-- d3441d
	sted3441d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3441d,
			Enable=>Enabled3441d,
			match=>matchd3441d,
			run=>run);

	Enabled3441d <= matchd3440d;
	-- d3442d
	sted3442d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3442d,
			Enable=>Enabled3442d,
			match=>matchd3442d,
			run=>run);

	Enabled3442d <= matchd3442d OR matchd3441d;
	-- d3443d
	sted3443d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3443d,
			Enable=>Enabled3443d,
			match=>matchd3443d,
			run=>run);

	Enabled3443d <= matchd3442d;
	-- d3444d
	sted3444d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3444d,
			Enable=>Enabled3444d,
			match=>matchd3444d,
			run=>run);

	Enabled3444d <= matchd3443d;
	-- d3445d
	sted3445d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3445d,
			Enable=>Enabled3445d,
			match=>matchd3445d,
			run=>run);

	Enabled3445d <= matchd3444d;
	-- d3446d
	sted3446d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3446d,
			Enable=>Enabled3446d,
			match=>matchd3446d,
			run=>run);

	reports(184) <= matchd3446d;
	Enabled3446d <= matchd3445d;
	-- d3447d
	sted3447d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3447d,
			Enable=>Enabled3447d,
			match=>matchd3447d,
			run=>run);

	-- d3448d
	sted3448d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3448d,
			Enable=>Enabled3448d,
			match=>matchd3448d,
			run=>run);

	Enabled3448d <= matchd3448d OR matchd3447d;
	-- d3449d
	sted3449d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3449d,
			Enable=>Enabled3449d,
			match=>matchd3449d,
			run=>run);

	Enabled3449d <= matchd3448d;
	-- d3450d
	sted3450d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3450d,
			Enable=>Enabled3450d,
			match=>matchd3450d,
			run=>run);

	Enabled3450d <= matchd3449d;
	-- d3451d
	sted3451d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3451d,
			Enable=>Enabled3451d,
			match=>matchd3451d,
			run=>run);

	Enabled3451d <= matchd3450d;
	-- d3452d
	sted3452d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3452d,
			Enable=>Enabled3452d,
			match=>matchd3452d,
			run=>run);

	Enabled3452d <= matchd3451d;
	-- d3453d
	sted3453d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3453d,
			Enable=>Enabled3453d,
			match=>matchd3453d,
			run=>run);

	Enabled3453d <= matchd3452d OR matchd3453d;
	-- d3454d
	sted3454d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3454d,
			Enable=>Enabled3454d,
			match=>matchd3454d,
			run=>run);

	Enabled3454d <= matchd3453d;
	-- d3455d
	sted3455d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3455d,
			Enable=>Enabled3455d,
			match=>matchd3455d,
			run=>run);

	Enabled3455d <= matchd3454d;
	-- d3456d
	sted3456d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3456d,
			Enable=>Enabled3456d,
			match=>matchd3456d,
			run=>run);

	Enabled3456d <= matchd3455d;
	-- d3457d
	sted3457d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3457d,
			Enable=>Enabled3457d,
			match=>matchd3457d,
			run=>run);

	reports(185) <= matchd3457d;
	Enabled3457d <= matchd3456d;
	-- d3458d
	sted3458d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3458d,
			Enable=>Enabled3458d,
			match=>matchd3458d,
			run=>run);

	-- d3459d
	sted3459d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3459d,
			Enable=>Enabled3459d,
			match=>matchd3459d,
			run=>run);

	Enabled3459d <= matchd3458d OR matchd3459d;
	-- d3460d
	sted3460d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3460d,
			Enable=>Enabled3460d,
			match=>matchd3460d,
			run=>run);

	Enabled3460d <= matchd3459d;
	-- d3461d
	sted3461d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3461d,
			Enable=>Enabled3461d,
			match=>matchd3461d,
			run=>run);

	Enabled3461d <= matchd3460d;
	-- d3462d
	sted3462d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3462d,
			Enable=>Enabled3462d,
			match=>matchd3462d,
			run=>run);

	Enabled3462d <= matchd3461d;
	-- d3463d
	sted3463d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3463d,
			Enable=>Enabled3463d,
			match=>matchd3463d,
			run=>run);

	Enabled3463d <= matchd3462d;
	-- d3464d
	sted3464d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3464d,
			Enable=>Enabled3464d,
			match=>matchd3464d,
			run=>run);

	Enabled3464d <= matchd3463d;
	-- d3465d
	sted3465d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3465d,
			Enable=>Enabled3465d,
			match=>matchd3465d,
			run=>run);

	Enabled3465d <= matchd3465d OR matchd3464d;
	-- d3466d
	sted3466d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3466d,
			Enable=>Enabled3466d,
			match=>matchd3466d,
			run=>run);

	Enabled3466d <= matchd3465d;
	-- d3467d
	sted3467d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3467d,
			Enable=>Enabled3467d,
			match=>matchd3467d,
			run=>run);

	Enabled3467d <= matchd3466d;
	-- d3468d
	sted3468d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3468d,
			Enable=>Enabled3468d,
			match=>matchd3468d,
			run=>run);

	Enabled3468d <= matchd3467d;
	-- d3469d
	sted3469d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3469d,
			Enable=>Enabled3469d,
			match=>matchd3469d,
			run=>run);

	reports(186) <= matchd3469d;
	Enabled3469d <= matchd3468d;
	-- d3470d
	sted3470d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3470d,
			Enable=>Enabled3470d,
			match=>matchd3470d,
			run=>run);

	-- d3471d
	sted3471d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3471d,
			Enable=>Enabled3471d,
			match=>matchd3471d,
			run=>run);

	Enabled3471d <= matchd3470d OR matchd3471d;
	-- d3472d
	sted3472d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3472d,
			Enable=>Enabled3472d,
			match=>matchd3472d,
			run=>run);

	Enabled3472d <= matchd3471d;
	-- d3473d
	sted3473d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3473d,
			Enable=>Enabled3473d,
			match=>matchd3473d,
			run=>run);

	Enabled3473d <= matchd3472d;
	-- d3474d
	sted3474d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3474d,
			Enable=>Enabled3474d,
			match=>matchd3474d,
			run=>run);

	Enabled3474d <= matchd3473d;
	-- d3475d
	sted3475d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3475d,
			Enable=>Enabled3475d,
			match=>matchd3475d,
			run=>run);

	Enabled3475d <= matchd3474d;
	-- d3476d
	sted3476d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3476d,
			Enable=>Enabled3476d,
			match=>matchd3476d,
			run=>run);

	Enabled3476d <= matchd3476d OR matchd3475d;
	-- d3477d
	sted3477d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3477d,
			Enable=>Enabled3477d,
			match=>matchd3477d,
			run=>run);

	Enabled3477d <= matchd3476d;
	-- d3478d
	sted3478d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3478d,
			Enable=>Enabled3478d,
			match=>matchd3478d,
			run=>run);

	Enabled3478d <= matchd3477d;
	-- d3479d
	sted3479d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3479d,
			Enable=>Enabled3479d,
			match=>matchd3479d,
			run=>run);

	Enabled3479d <= matchd3478d;
	-- d3480d
	sted3480d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3480d,
			Enable=>Enabled3480d,
			match=>matchd3480d,
			run=>run);

	Enabled3480d <= matchd3479d;
	-- d3481d
	sted3481d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3481d,
			Enable=>Enabled3481d,
			match=>matchd3481d,
			run=>run);

	Enabled3481d <= matchd3481d OR matchd3480d;
	-- d3482d
	sted3482d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3482d,
			Enable=>Enabled3482d,
			match=>matchd3482d,
			run=>run);

	Enabled3482d <= matchd3481d;
	-- d3483d
	sted3483d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3483d,
			Enable=>Enabled3483d,
			match=>matchd3483d,
			run=>run);

	Enabled3483d <= matchd3482d;
	-- d3484d
	sted3484d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3484d,
			Enable=>Enabled3484d,
			match=>matchd3484d,
			run=>run);

	Enabled3484d <= matchd3483d;
	-- d3485d
	sted3485d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3485d,
			Enable=>Enabled3485d,
			match=>matchd3485d,
			run=>run);

	reports(187) <= matchd3485d;
	Enabled3485d <= matchd3484d;
	-- d3486d
	sted3486d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3486d,
			Enable=>Enabled3486d,
			match=>matchd3486d,
			run=>run);

	-- d3487d
	sted3487d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3487d,
			Enable=>Enabled3487d,
			match=>matchd3487d,
			run=>run);

	Enabled3487d <= matchd3487d OR matchd3486d;
	-- d3488d
	sted3488d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3488d,
			Enable=>Enabled3488d,
			match=>matchd3488d,
			run=>run);

	Enabled3488d <= matchd3487d;
	-- d3489d
	sted3489d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3489d,
			Enable=>Enabled3489d,
			match=>matchd3489d,
			run=>run);

	Enabled3489d <= matchd3488d;
	-- d3490d
	sted3490d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3490d,
			Enable=>Enabled3490d,
			match=>matchd3490d,
			run=>run);

	Enabled3490d <= matchd3489d;
	-- d3491d
	sted3491d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3491d,
			Enable=>Enabled3491d,
			match=>matchd3491d,
			run=>run);

	Enabled3491d <= matchd3490d;
	-- d3492d
	sted3492d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3492d,
			Enable=>Enabled3492d,
			match=>matchd3492d,
			run=>run);

	Enabled3492d <= matchd3491d;
	-- d3493d
	sted3493d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3493d,
			Enable=>Enabled3493d,
			match=>matchd3493d,
			run=>run);

	Enabled3493d <= matchd3492d OR matchd3493d;
	-- d3494d
	sted3494d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3494d,
			Enable=>Enabled3494d,
			match=>matchd3494d,
			run=>run);

	Enabled3494d <= matchd3493d;
	-- d3495d
	sted3495d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3495d,
			Enable=>Enabled3495d,
			match=>matchd3495d,
			run=>run);

	Enabled3495d <= matchd3494d;
	-- d3496d
	sted3496d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3496d,
			Enable=>Enabled3496d,
			match=>matchd3496d,
			run=>run);

	Enabled3496d <= matchd3495d;
	-- d3497d
	sted3497d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3497d,
			Enable=>Enabled3497d,
			match=>matchd3497d,
			run=>run);

	Enabled3497d <= matchd3496d;
	-- d3498d
	sted3498d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3498d,
			Enable=>Enabled3498d,
			match=>matchd3498d,
			run=>run);

	Enabled3498d <= matchd3498d OR matchd3497d;
	-- d3499d
	sted3499d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3499d,
			Enable=>Enabled3499d,
			match=>matchd3499d,
			run=>run);

	Enabled3499d <= matchd3498d;
	-- d3500d
	sted3500d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3500d,
			Enable=>Enabled3500d,
			match=>matchd3500d,
			run=>run);

	Enabled3500d <= matchd3499d;
	-- d3501d
	sted3501d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3501d,
			Enable=>Enabled3501d,
			match=>matchd3501d,
			run=>run);

	Enabled3501d <= matchd3500d;
	-- d3502d
	sted3502d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3502d,
			Enable=>Enabled3502d,
			match=>matchd3502d,
			run=>run);

	reports(188) <= matchd3502d;
	Enabled3502d <= matchd3501d;
	-- d3503d
	sted3503d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3503d,
			Enable=>Enabled3503d,
			match=>matchd3503d,
			run=>run);

	-- d3504d
	sted3504d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3504d,
			Enable=>Enabled3504d,
			match=>matchd3504d,
			run=>run);

	Enabled3504d <= matchd3503d;
	-- d3505d
	sted3505d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3505d,
			Enable=>Enabled3505d,
			match=>matchd3505d,
			run=>run);

	Enabled3505d <= matchd3504d;
	-- d3506d
	sted3506d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3506d,
			Enable=>Enabled3506d,
			match=>matchd3506d,
			run=>run);

	Enabled3506d <= matchd3505d;
	-- d3507d
	sted3507d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3507d,
			Enable=>Enabled3507d,
			match=>matchd3507d,
			run=>run);

	Enabled3507d <= matchd3506d;
	-- d3508d
	sted3508d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3508d,
			Enable=>Enabled3508d,
			match=>matchd3508d,
			run=>run);

	Enabled3508d <= matchd3507d;
	-- d3509d
	sted3509d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3509d,
			Enable=>Enabled3509d,
			match=>matchd3509d,
			run=>run);

	Enabled3509d <= matchd3508d;
	-- d3510d
	sted3510d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3510d,
			Enable=>Enabled3510d,
			match=>matchd3510d,
			run=>run);

	Enabled3510d <= matchd3509d;
	-- d3511d
	sted3511d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3511d,
			Enable=>Enabled3511d,
			match=>matchd3511d,
			run=>run);

	Enabled3511d <= matchd3510d;
	-- d3512d
	sted3512d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3512d,
			Enable=>Enabled3512d,
			match=>matchd3512d,
			run=>run);

	Enabled3512d <= matchd3511d;
	-- d3513d
	sted3513d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3513d,
			Enable=>Enabled3513d,
			match=>matchd3513d,
			run=>run);

	Enabled3513d <= matchd3512d;
	-- d3514d
	sted3514d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3514d,
			Enable=>Enabled3514d,
			match=>matchd3514d,
			run=>run);

	Enabled3514d <= matchd3513d;
	-- d3515d
	sted3515d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3515d,
			Enable=>Enabled3515d,
			match=>matchd3515d,
			run=>run);

	Enabled3515d <= matchd3515d OR matchd3514d;
	-- d3516d
	sted3516d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3516d,
			Enable=>Enabled3516d,
			match=>matchd3516d,
			run=>run);

	Enabled3516d <= matchd3515d;
	-- d3517d
	sted3517d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3517d,
			Enable=>Enabled3517d,
			match=>matchd3517d,
			run=>run);

	Enabled3517d <= matchd3516d;
	-- d3518d
	sted3518d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3518d,
			Enable=>Enabled3518d,
			match=>matchd3518d,
			run=>run);

	Enabled3518d <= matchd3517d;
	-- d3519d
	sted3519d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3519d,
			Enable=>Enabled3519d,
			match=>matchd3519d,
			run=>run);

	reports(189) <= matchd3519d;
	Enabled3519d <= matchd3518d;
	-- d3520d
	sted3520d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3520d,
			Enable=>Enabled3520d,
			match=>matchd3520d,
			run=>run);

	-- d3521d
	sted3521d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3521d,
			Enable=>Enabled3521d,
			match=>matchd3521d,
			run=>run);

	Enabled3521d <= matchd3521d OR matchd3520d;
	-- d3522d
	sted3522d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3522d,
			Enable=>Enabled3522d,
			match=>matchd3522d,
			run=>run);

	Enabled3522d <= matchd3521d;
	-- d3523d
	sted3523d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3523d,
			Enable=>Enabled3523d,
			match=>matchd3523d,
			run=>run);

	Enabled3523d <= matchd3522d;
	-- d3524d
	sted3524d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3524d,
			Enable=>Enabled3524d,
			match=>matchd3524d,
			run=>run);

	Enabled3524d <= matchd3523d;
	-- d3525d
	sted3525d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3525d,
			Enable=>Enabled3525d,
			match=>matchd3525d,
			run=>run);

	Enabled3525d <= matchd3524d;
	-- d3526d
	sted3526d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3526d,
			Enable=>Enabled3526d,
			match=>matchd3526d,
			run=>run);

	Enabled3526d <= matchd3525d;
	-- d3527d
	sted3527d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3527d,
			Enable=>Enabled3527d,
			match=>matchd3527d,
			run=>run);

	Enabled3527d <= matchd3526d;
	-- d3528d
	sted3528d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3528d,
			Enable=>Enabled3528d,
			match=>matchd3528d,
			run=>run);

	Enabled3528d <= matchd3527d;
	-- d3529d
	sted3529d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3529d,
			Enable=>Enabled3529d,
			match=>matchd3529d,
			run=>run);

	Enabled3529d <= matchd3528d;
	-- d3530d
	sted3530d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3530d,
			Enable=>Enabled3530d,
			match=>matchd3530d,
			run=>run);

	Enabled3530d <= matchd3529d OR matchd3530d;
	-- d3531d
	sted3531d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3531d,
			Enable=>Enabled3531d,
			match=>matchd3531d,
			run=>run);

	Enabled3531d <= matchd3530d;
	-- d3532d
	sted3532d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3532d,
			Enable=>Enabled3532d,
			match=>matchd3532d,
			run=>run);

	Enabled3532d <= matchd3531d;
	-- d3533d
	sted3533d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3533d,
			Enable=>Enabled3533d,
			match=>matchd3533d,
			run=>run);

	Enabled3533d <= matchd3532d;
	-- d3534d
	sted3534d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3534d,
			Enable=>Enabled3534d,
			match=>matchd3534d,
			run=>run);

	Enabled3534d <= matchd3533d;
	-- d3535d
	sted3535d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3535d,
			Enable=>Enabled3535d,
			match=>matchd3535d,
			run=>run);

	Enabled3535d <= matchd3534d;
	-- d3536d
	sted3536d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3536d,
			Enable=>Enabled3536d,
			match=>matchd3536d,
			run=>run);

	Enabled3536d <= matchd3536d OR matchd3535d;
	-- d3537d
	sted3537d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3537d,
			Enable=>Enabled3537d,
			match=>matchd3537d,
			run=>run);

	Enabled3537d <= matchd3536d;
	-- d3538d
	sted3538d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3538d,
			Enable=>Enabled3538d,
			match=>matchd3538d,
			run=>run);

	Enabled3538d <= matchd3537d;
	-- d3539d
	sted3539d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3539d,
			Enable=>Enabled3539d,
			match=>matchd3539d,
			run=>run);

	Enabled3539d <= matchd3538d;
	-- d3540d
	sted3540d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3540d,
			Enable=>Enabled3540d,
			match=>matchd3540d,
			run=>run);

	Enabled3540d <= matchd3539d;
	-- d3541d
	sted3541d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3541d,
			Enable=>Enabled3541d,
			match=>matchd3541d,
			run=>run);

	reports(190) <= matchd3541d;
	Enabled3541d <= matchd3540d;
	-- d3542d
	sted3542d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3542d,
			Enable=>Enabled3542d,
			match=>matchd3542d,
			run=>run);

	-- d3543d
	sted3543d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3543d,
			Enable=>Enabled3543d,
			match=>matchd3543d,
			run=>run);

	Enabled3543d <= matchd3542d OR matchd3543d;
	-- d3544d
	sted3544d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3544d,
			Enable=>Enabled3544d,
			match=>matchd3544d,
			run=>run);

	Enabled3544d <= matchd3543d;
	-- d3545d
	sted3545d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3545d,
			Enable=>Enabled3545d,
			match=>matchd3545d,
			run=>run);

	Enabled3545d <= matchd3544d;
	-- d3546d
	sted3546d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3546d,
			Enable=>Enabled3546d,
			match=>matchd3546d,
			run=>run);

	Enabled3546d <= matchd3545d;
	-- d3547d
	sted3547d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3547d,
			Enable=>Enabled3547d,
			match=>matchd3547d,
			run=>run);

	Enabled3547d <= matchd3546d;
	-- d3548d
	sted3548d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3548d,
			Enable=>Enabled3548d,
			match=>matchd3548d,
			run=>run);

	Enabled3548d <= matchd3547d OR matchd3548d;
	-- d3549d
	sted3549d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3549d,
			Enable=>Enabled3549d,
			match=>matchd3549d,
			run=>run);

	Enabled3549d <= matchd3548d;
	-- d3550d
	sted3550d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3550d,
			Enable=>Enabled3550d,
			match=>matchd3550d,
			run=>run);

	Enabled3550d <= matchd3549d;
	-- d3551d
	sted3551d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3551d,
			Enable=>Enabled3551d,
			match=>matchd3551d,
			run=>run);

	Enabled3551d <= matchd3550d;
	-- d3552d
	sted3552d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3552d,
			Enable=>Enabled3552d,
			match=>matchd3552d,
			run=>run);

	Enabled3552d <= matchd3551d;
	-- d3553d
	sted3553d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3553d,
			Enable=>Enabled3553d,
			match=>matchd3553d,
			run=>run);

	Enabled3553d <= matchd3553d OR matchd3552d;
	-- d3554d
	sted3554d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3554d,
			Enable=>Enabled3554d,
			match=>matchd3554d,
			run=>run);

	Enabled3554d <= matchd3553d;
	-- d3555d
	sted3555d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3555d,
			Enable=>Enabled3555d,
			match=>matchd3555d,
			run=>run);

	Enabled3555d <= matchd3554d;
	-- d3556d
	sted3556d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3556d,
			Enable=>Enabled3556d,
			match=>matchd3556d,
			run=>run);

	Enabled3556d <= matchd3555d;
	-- d3557d
	sted3557d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3557d,
			Enable=>Enabled3557d,
			match=>matchd3557d,
			run=>run);

	reports(191) <= matchd3557d;
	Enabled3557d <= matchd3556d;
	-- d3558d
	sted3558d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3558d,
			Enable=>Enabled3558d,
			match=>matchd3558d,
			run=>run);

	-- d3559d
	sted3559d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3559d,
			Enable=>Enabled3559d,
			match=>matchd3559d,
			run=>run);

	Enabled3559d <= matchd3558d OR matchd3559d;
	-- d3560d
	sted3560d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3560d,
			Enable=>Enabled3560d,
			match=>matchd3560d,
			run=>run);

	Enabled3560d <= matchd3559d;
	-- d3561d
	sted3561d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3561d,
			Enable=>Enabled3561d,
			match=>matchd3561d,
			run=>run);

	Enabled3561d <= matchd3560d;
	-- d3562d
	sted3562d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3562d,
			Enable=>Enabled3562d,
			match=>matchd3562d,
			run=>run);

	Enabled3562d <= matchd3561d;
	-- d3563d
	sted3563d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3563d,
			Enable=>Enabled3563d,
			match=>matchd3563d,
			run=>run);

	Enabled3563d <= matchd3562d;
	-- d3564d
	sted3564d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3564d,
			Enable=>Enabled3564d,
			match=>matchd3564d,
			run=>run);

	Enabled3564d <= matchd3563d;
	-- d3565d
	sted3565d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3565d,
			Enable=>Enabled3565d,
			match=>matchd3565d,
			run=>run);

	Enabled3565d <= matchd3564d OR matchd3565d;
	-- d3566d
	sted3566d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3566d,
			Enable=>Enabled3566d,
			match=>matchd3566d,
			run=>run);

	Enabled3566d <= matchd3565d;
	-- d3567d
	sted3567d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3567d,
			Enable=>Enabled3567d,
			match=>matchd3567d,
			run=>run);

	Enabled3567d <= matchd3566d;
	-- d3568d
	sted3568d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3568d,
			Enable=>Enabled3568d,
			match=>matchd3568d,
			run=>run);

	Enabled3568d <= matchd3567d;
	-- d3569d
	sted3569d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3569d,
			Enable=>Enabled3569d,
			match=>matchd3569d,
			run=>run);

	Enabled3569d <= matchd3568d;
	-- d3570d
	sted3570d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3570d,
			Enable=>Enabled3570d,
			match=>matchd3570d,
			run=>run);

	Enabled3570d <= matchd3569d;
	-- d3571d
	sted3571d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3571d,
			Enable=>Enabled3571d,
			match=>matchd3571d,
			run=>run);

	Enabled3571d <= matchd3571d OR matchd3570d;
	-- d3572d
	sted3572d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3572d,
			Enable=>Enabled3572d,
			match=>matchd3572d,
			run=>run);

	Enabled3572d <= matchd3571d;
	-- d3573d
	sted3573d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3573d,
			Enable=>Enabled3573d,
			match=>matchd3573d,
			run=>run);

	Enabled3573d <= matchd3572d;
	-- d3574d
	sted3574d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3574d,
			Enable=>Enabled3574d,
			match=>matchd3574d,
			run=>run);

	Enabled3574d <= matchd3573d;
	-- d3575d
	sted3575d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3575d,
			Enable=>Enabled3575d,
			match=>matchd3575d,
			run=>run);

	Enabled3575d <= matchd3574d;
	-- d3576d
	sted3576d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3576d,
			Enable=>Enabled3576d,
			match=>matchd3576d,
			run=>run);

	Enabled3576d <= matchd3575d;
	-- d3577d
	sted3577d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3577d,
			Enable=>Enabled3577d,
			match=>matchd3577d,
			run=>run);

	reports(192) <= matchd3577d;
	Enabled3577d <= matchd3576d;
	-- d3578d
	sted3578d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3578d,
			Enable=>Enabled3578d,
			match=>matchd3578d,
			run=>run);

	-- d3579d
	sted3579d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3579d,
			Enable=>Enabled3579d,
			match=>matchd3579d,
			run=>run);

	Enabled3579d <= matchd3579d OR matchd3578d;
	-- d3580d
	sted3580d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3580d,
			Enable=>Enabled3580d,
			match=>matchd3580d,
			run=>run);

	Enabled3580d <= matchd3579d;
	-- d3581d
	sted3581d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3581d,
			Enable=>Enabled3581d,
			match=>matchd3581d,
			run=>run);

	Enabled3581d <= matchd3580d;
	-- d3582d
	sted3582d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3582d,
			Enable=>Enabled3582d,
			match=>matchd3582d,
			run=>run);

	Enabled3582d <= matchd3581d;
	-- d3583d
	sted3583d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3583d,
			Enable=>Enabled3583d,
			match=>matchd3583d,
			run=>run);

	Enabled3583d <= matchd3582d;
	-- d3584d
	sted3584d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3584d,
			Enable=>Enabled3584d,
			match=>matchd3584d,
			run=>run);

	Enabled3584d <= matchd3583d OR matchd3584d;
	-- d3585d
	sted3585d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3585d,
			Enable=>Enabled3585d,
			match=>matchd3585d,
			run=>run);

	Enabled3585d <= matchd3584d;
	-- d3586d
	sted3586d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3586d,
			Enable=>Enabled3586d,
			match=>matchd3586d,
			run=>run);

	Enabled3586d <= matchd3585d;
	-- d3587d
	sted3587d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3587d,
			Enable=>Enabled3587d,
			match=>matchd3587d,
			run=>run);

	Enabled3587d <= matchd3586d;
	-- d3588d
	sted3588d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3588d,
			Enable=>Enabled3588d,
			match=>matchd3588d,
			run=>run);

	Enabled3588d <= matchd3587d;
	-- d3589d
	sted3589d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3589d,
			Enable=>Enabled3589d,
			match=>matchd3589d,
			run=>run);

	Enabled3589d <= matchd3588d OR matchd3589d;
	-- d3590d
	sted3590d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3590d,
			Enable=>Enabled3590d,
			match=>matchd3590d,
			run=>run);

	Enabled3590d <= matchd3589d;
	-- d3591d
	sted3591d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3591d,
			Enable=>Enabled3591d,
			match=>matchd3591d,
			run=>run);

	Enabled3591d <= matchd3590d;
	-- d3592d
	sted3592d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3592d,
			Enable=>Enabled3592d,
			match=>matchd3592d,
			run=>run);

	Enabled3592d <= matchd3591d;
	-- d3593d
	sted3593d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3593d,
			Enable=>Enabled3593d,
			match=>matchd3593d,
			run=>run);

	Enabled3593d <= matchd3592d;
	-- d3594d
	sted3594d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3594d,
			Enable=>Enabled3594d,
			match=>matchd3594d,
			run=>run);

	reports(193) <= matchd3594d;
	Enabled3594d <= matchd3593d;
	-- d3595d
	sted3595d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3595d,
			Enable=>Enabled3595d,
			match=>matchd3595d,
			run=>run);

	-- d3596d
	sted3596d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3596d,
			Enable=>Enabled3596d,
			match=>matchd3596d,
			run=>run);

	Enabled3596d <= matchd3596d OR matchd3595d;
	-- d3597d
	sted3597d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3597d,
			Enable=>Enabled3597d,
			match=>matchd3597d,
			run=>run);

	Enabled3597d <= matchd3596d;
	-- d3598d
	sted3598d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3598d,
			Enable=>Enabled3598d,
			match=>matchd3598d,
			run=>run);

	Enabled3598d <= matchd3597d;
	-- d3599d
	sted3599d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3599d,
			Enable=>Enabled3599d,
			match=>matchd3599d,
			run=>run);

	Enabled3599d <= matchd3598d;
	-- d3600d
	sted3600d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3600d,
			Enable=>Enabled3600d,
			match=>matchd3600d,
			run=>run);

	Enabled3600d <= matchd3599d;
	-- d3601d
	sted3601d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3601d,
			Enable=>Enabled3601d,
			match=>matchd3601d,
			run=>run);

	Enabled3601d <= matchd3601d OR matchd3600d;
	-- d3602d
	sted3602d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3602d,
			Enable=>Enabled3602d,
			match=>matchd3602d,
			run=>run);

	Enabled3602d <= matchd3601d;
	-- d3603d
	sted3603d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3603d,
			Enable=>Enabled3603d,
			match=>matchd3603d,
			run=>run);

	Enabled3603d <= matchd3602d;
	-- d3604d
	sted3604d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3604d,
			Enable=>Enabled3604d,
			match=>matchd3604d,
			run=>run);

	Enabled3604d <= matchd3603d;
	-- d3605d
	sted3605d : ste_sim
	port map(char_in=>data_in,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectord3605d,
			Enable=>Enabled3605d,
			match=>matchd3605d,
			run=>run);

	reports(194) <= matchd3605d;
	Enabled3605d <= matchd3604d;
	

	-- reset_n <= not reset;--VINH commented this since it seems reset_n will not be used

	
	--- ORs
	-- d269d
	matchd269d <= matchd251d OR matchd268d;
	reports(195) <= matchd269d;
	
	-- d313d
	matchd313d <= matchd312d OR matchd297d;
	reports(196) <= matchd313d;
	
	-- d356d
	matchd356d <= matchd340d OR matchd355d;
	reports(197) <= matchd356d;
	
	-- d433d
	matchd433d <= matchd390d OR matchd411d OR matchd432d;
	reports(198) <= matchd433d;
	
	-- d505d
	matchd505d <= matchd484d OR matchd504d OR matchd464d;
	reports(199) <= matchd505d;
	
	-- d554d
	matchd554d <= matchd553d OR matchd537d;
	reports(200) <= matchd554d;
	
	-- d626d
	matchd626d <= matchd605d OR matchd585d OR matchd625d;
	reports(201) <= matchd626d;
	
	-- d725d
	matchd725d <= matchd707d OR matchd724d;
	reports(202) <= matchd725d;
	
	-- d818d
	matchd818d <= matchd802d OR matchd817d;
	reports(203) <= matchd818d;
	
	-- d906d
	matchd906d <= matchd905d OR matchd863d OR matchd884d;
	reports(204) <= matchd906d;
	
	-- d985d
	matchd985d <= matchd970d OR matchd984d;
	reports(205) <= matchd985d;
	
	-- d1119d
	matchd1119d <= matchd1118d OR matchd1101d;
	reports(206) <= matchd1119d;
	
	-- d1299d
	matchd1299d <= matchd1298d OR matchd1282d;
	reports(207) <= matchd1299d;
	
	-- d1763d
	matchd1763d <= matchd1762d OR matchd1745d;
	reports(208) <= matchd1763d;
	
	-- d1851d
	matchd1851d <= matchd1850d OR matchd1832d OR matchd1814d;
	reports(209) <= matchd1851d;
	
	-- d2324d
	matchd2324d <= matchd2323d OR matchd2307d;
	reports(210) <= matchd2324d;
	
	-- d2397d
	matchd2397d <= matchd2396d OR matchd2381d;
	reports(211) <= matchd2397d;
	
	-- d2836d
	matchd2836d <= matchd2835d OR matchd2818d;
	reports(212) <= matchd2836d;
	
	-- d2869d
	matchd2869d <= matchd2868d OR matchd2852d;
	reports(213) <= matchd2869d;
	
	-- d3058d
	matchd3058d <= matchd3040d OR matchd3057d;
	reports(214) <= matchd3058d;
	
	-- d3116d
	matchd3116d <= matchd3077d OR matchd3115d OR matchd3096d;
	reports(215) <= matchd3116d;
	
	-- d3182d
	matchd3182d <= matchd3165d OR matchd3181d;
	reports(216) <= matchd3182d;
	
	-- d3295d
	matchd3295d <= matchd3277d OR matchd3294d;
	reports(217) <= matchd3295d;
	
	
	--- ANDs
	--- Counters
end Structure;